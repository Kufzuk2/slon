module tile_rom (                       //невскрытая клетка
  input  wire    [13:0]     addr,
  output wire    [11:0]     word
);

  logic [11:0] rom [(25 * 25)];

  assign word = rom[addr];

  initial begin
rom[0] = 12'hfff
rom[1] = 12'hfff
rom[2] = 12'hfff
rom[3] = 12'hfff
rom[4] = 12'hfff
rom[5] = 12'hfff
rom[6] = 12'hfff
rom[7] = 12'hfff
rom[8] = 12'hfff
rom[9] = 12'hfff
rom[10] = 12'hfff
rom[11] = 12'hfff
rom[12] = 12'hfff
rom[13] = 12'hfff
rom[14] = 12'hfff
rom[15] = 12'hfff
rom[16] = 12'hfff
rom[17] = 12'hfff
rom[18] = 12'hfff
rom[19] = 12'hfff
rom[20] = 12'hfff
rom[21] = 12'hfff
rom[22] = 12'hfff
rom[23] = 12'hfff
rom[24] = 12'h777
rom[25] = 12'hfff
rom[26] = 12'hfff
rom[27] = 12'hfff
rom[28] = 12'hfff
rom[29] = 12'hfff
rom[30] = 12'hfff
rom[31] = 12'hfff
rom[32] = 12'hfff
rom[33] = 12'hfff
rom[34] = 12'hfff
rom[35] = 12'hfff
rom[36] = 12'hfff
rom[37] = 12'hfff
rom[38] = 12'hfff
rom[39] = 12'hfff
rom[40] = 12'hfff
rom[41] = 12'hfff
rom[42] = 12'hfff
rom[43] = 12'hfff
rom[44] = 12'hfff
rom[45] = 12'hfff
rom[46] = 12'hfff
rom[47] = 12'hfff
rom[48] = 12'h777
rom[49] = 12'h777
rom[50] = 12'hfff
rom[51] = 12'hfff
rom[52] = 12'hfff
rom[53] = 12'hfff
rom[54] = 12'hfff
rom[55] = 12'hfff
rom[56] = 12'hfff
rom[57] = 12'hfff
rom[58] = 12'hfff
rom[59] = 12'hfff
rom[60] = 12'hfff
rom[61] = 12'hfff
rom[62] = 12'hfff
rom[63] = 12'hfff
rom[64] = 12'hfff
rom[65] = 12'hfff
rom[66] = 12'hfff
rom[67] = 12'hfff
rom[68] = 12'hfff
rom[69] = 12'hfff
rom[70] = 12'hfff
rom[71] = 12'hfff
rom[72] = 12'h777
rom[73] = 12'h777
rom[74] = 12'h777
rom[75] = 12'hfff
rom[76] = 12'hfff
rom[77] = 12'hfff
rom[78] = 12'hccc
rom[79] = 12'hccc
rom[80] = 12'hccc
rom[81] = 12'hccc
rom[82] = 12'hccc
rom[83] = 12'hccc
rom[84] = 12'hccc
rom[85] = 12'hccc
rom[86] = 12'hccc
rom[87] = 12'hccc
rom[88] = 12'hccc
rom[89] = 12'hccc
rom[90] = 12'hccc
rom[91] = 12'hccc
rom[92] = 12'hccc
rom[93] = 12'hccc
rom[94] = 12'hccc
rom[95] = 12'hccc
rom[96] = 12'h777
rom[97] = 12'h777
rom[98] = 12'h777
rom[99] = 12'h777
rom[100] = 12'hfff
rom[101] = 12'hfff
rom[102] = 12'hfff
rom[103] = 12'hccc
rom[104] = 12'hccc
rom[105] = 12'hccc
rom[106] = 12'hccc
rom[107] = 12'hccc
rom[108] = 12'hccc
rom[109] = 12'hccc
rom[110] = 12'hccc
rom[111] = 12'hccc
rom[112] = 12'hccc
rom[113] = 12'hccc
rom[114] = 12'hccc
rom[115] = 12'hccc
rom[116] = 12'hccc
rom[117] = 12'hccc
rom[118] = 12'hccc
rom[119] = 12'hccc
rom[120] = 12'hccc
rom[121] = 12'h777
rom[122] = 12'h777
rom[123] = 12'h777
rom[124] = 12'h777
rom[125] = 12'hfff
rom[126] = 12'hfff
rom[127] = 12'hfff
rom[128] = 12'hccc
rom[129] = 12'hccc
rom[130] = 12'hccc
rom[131] = 12'hccc
rom[132] = 12'hccc
rom[133] = 12'hccc
rom[134] = 12'hccc
rom[135] = 12'hccc
rom[136] = 12'hccc
rom[137] = 12'hccc
rom[138] = 12'hccc
rom[139] = 12'hccc
rom[140] = 12'hccc
rom[141] = 12'hccc
rom[142] = 12'hccc
rom[143] = 12'hccc
rom[144] = 12'hccc
rom[145] = 12'hccc
rom[146] = 12'h777
rom[147] = 12'h777
rom[148] = 12'h777
rom[149] = 12'h777
rom[150] = 12'hfff
rom[151] = 12'hfff
rom[152] = 12'hfff
rom[153] = 12'hccc
rom[154] = 12'hccc
rom[155] = 12'hccc
rom[156] = 12'hccc
rom[157] = 12'hccc
rom[158] = 12'hccc
rom[159] = 12'hccc
rom[160] = 12'hccc
rom[161] = 12'hccc
rom[162] = 12'hccc
rom[163] = 12'hccc
rom[164] = 12'hccc
rom[165] = 12'hccc
rom[166] = 12'hccc
rom[167] = 12'hccc
rom[168] = 12'hccc
rom[169] = 12'hccc
rom[170] = 12'hccc
rom[171] = 12'h777
rom[172] = 12'h777
rom[173] = 12'h777
rom[174] = 12'h777
rom[175] = 12'hfff
rom[176] = 12'hfff
rom[177] = 12'hfff
rom[178] = 12'hccc
rom[179] = 12'hccc
rom[180] = 12'hccc
rom[181] = 12'hccc
rom[182] = 12'hccc
rom[183] = 12'hccc
rom[184] = 12'hccc
rom[185] = 12'hccc
rom[186] = 12'hccc
rom[187] = 12'hccc
rom[188] = 12'hccc
rom[189] = 12'hccc
rom[190] = 12'hccc
rom[191] = 12'hccc
rom[192] = 12'hccc
rom[193] = 12'hccc
rom[194] = 12'hccc
rom[195] = 12'hccc
rom[196] = 12'h777
rom[197] = 12'h777
rom[198] = 12'h777
rom[199] = 12'h777
rom[200] = 12'hfff
rom[201] = 12'hfff
rom[202] = 12'hfff
rom[203] = 12'hccc
rom[204] = 12'hccc
rom[205] = 12'hccc
rom[206] = 12'hccc
rom[207] = 12'hccc
rom[208] = 12'hccc
rom[209] = 12'hccc
rom[210] = 12'hccc
rom[211] = 12'hccc
rom[212] = 12'hccc
rom[213] = 12'hccc
rom[214] = 12'hccc
rom[215] = 12'hccc
rom[216] = 12'hccc
rom[217] = 12'hccc
rom[218] = 12'hccc
rom[219] = 12'hccc
rom[220] = 12'hccc
rom[221] = 12'h777
rom[222] = 12'h777
rom[223] = 12'h777
rom[224] = 12'h777
rom[225] = 12'hfff
rom[226] = 12'hfff
rom[227] = 12'hfff
rom[228] = 12'hccc
rom[229] = 12'hccc
rom[230] = 12'hccc
rom[231] = 12'hccc
rom[232] = 12'hccc
rom[233] = 12'hccc
rom[234] = 12'hccc
rom[235] = 12'hccc
rom[236] = 12'hccc
rom[237] = 12'hccc
rom[238] = 12'hccc
rom[239] = 12'hccc
rom[240] = 12'hccc
rom[241] = 12'hccc
rom[242] = 12'hccc
rom[243] = 12'hccc
rom[244] = 12'hccc
rom[245] = 12'hccc
rom[246] = 12'h777
rom[247] = 12'h777
rom[248] = 12'h777
rom[249] = 12'h777
rom[250] = 12'hfff
rom[251] = 12'hfff
rom[252] = 12'hfff
rom[253] = 12'hccc
rom[254] = 12'hccc
rom[255] = 12'hccc
rom[256] = 12'hccc
rom[257] = 12'hccc
rom[258] = 12'hccc
rom[259] = 12'hccc
rom[260] = 12'hccc
rom[261] = 12'hccc
rom[262] = 12'hccc
rom[263] = 12'hccc
rom[264] = 12'hccc
rom[265] = 12'hccc
rom[266] = 12'hccc
rom[267] = 12'hccc
rom[268] = 12'hccc
rom[269] = 12'hccc
rom[270] = 12'hccc
rom[271] = 12'h777
rom[272] = 12'h777
rom[273] = 12'h777
rom[274] = 12'h777
rom[275] = 12'hfff
rom[276] = 12'hfff
rom[277] = 12'hfff
rom[278] = 12'hccc
rom[279] = 12'hccc
rom[280] = 12'hccc
rom[281] = 12'hccc
rom[282] = 12'hccc
rom[283] = 12'hccc
rom[284] = 12'hccc
rom[285] = 12'hccc
rom[286] = 12'hccc
rom[287] = 12'hccc
rom[288] = 12'hccc
rom[289] = 12'hccc
rom[290] = 12'hccc
rom[291] = 12'hccc
rom[292] = 12'hccc
rom[293] = 12'hccc
rom[294] = 12'hccc
rom[295] = 12'hccc
rom[296] = 12'h777
rom[297] = 12'h777
rom[298] = 12'h777
rom[299] = 12'h777
rom[300] = 12'hfff
rom[301] = 12'hfff
rom[302] = 12'hfff
rom[303] = 12'hccc
rom[304] = 12'hccc
rom[305] = 12'hccc
rom[306] = 12'hccc
rom[307] = 12'hccc
rom[308] = 12'hccc
rom[309] = 12'hccc
rom[310] = 12'hccc
rom[311] = 12'hccc
rom[312] = 12'hccc
rom[313] = 12'hccc
rom[314] = 12'hccc
rom[315] = 12'hccc
rom[316] = 12'hccc
rom[317] = 12'hccc
rom[318] = 12'hccc
rom[319] = 12'hccc
rom[320] = 12'hccc
rom[321] = 12'h777
rom[322] = 12'h777
rom[323] = 12'h777
rom[324] = 12'h777
rom[325] = 12'hfff
rom[326] = 12'hfff
rom[327] = 12'hfff
rom[328] = 12'hccc
rom[329] = 12'hccc
rom[330] = 12'hccc
rom[331] = 12'hccc
rom[332] = 12'hccc
rom[333] = 12'hccc
rom[334] = 12'hccc
rom[335] = 12'hccc
rom[336] = 12'hccc
rom[337] = 12'hccc
rom[338] = 12'hccc
rom[339] = 12'hccc
rom[340] = 12'hccc
rom[341] = 12'hccc
rom[342] = 12'hccc
rom[343] = 12'hccc
rom[344] = 12'hccc
rom[345] = 12'hccc
rom[346] = 12'h777
rom[347] = 12'h777
rom[348] = 12'h777
rom[349] = 12'h777
rom[350] = 12'hfff
rom[351] = 12'hfff
rom[352] = 12'hfff
rom[353] = 12'hccc
rom[354] = 12'hccc
rom[355] = 12'hccc
rom[356] = 12'hccc
rom[357] = 12'hccc
rom[358] = 12'hccc
rom[359] = 12'hccc
rom[360] = 12'hccc
rom[361] = 12'hccc
rom[362] = 12'hccc
rom[363] = 12'hccc
rom[364] = 12'hccc
rom[365] = 12'hccc
rom[366] = 12'hccc
rom[367] = 12'hccc
rom[368] = 12'hccc
rom[369] = 12'hccc
rom[370] = 12'hccc
rom[371] = 12'h777
rom[372] = 12'h777
rom[373] = 12'h777
rom[374] = 12'h777
rom[375] = 12'hfff
rom[376] = 12'hfff
rom[377] = 12'hfff
rom[378] = 12'hccc
rom[379] = 12'hccc
rom[380] = 12'hccc
rom[381] = 12'hccc
rom[382] = 12'hccc
rom[383] = 12'hccc
rom[384] = 12'hccc
rom[385] = 12'hccc
rom[386] = 12'hccc
rom[387] = 12'hccc
rom[388] = 12'hccc
rom[389] = 12'hccc
rom[390] = 12'hccc
rom[391] = 12'hccc
rom[392] = 12'hccc
rom[393] = 12'hccc
rom[394] = 12'hccc
rom[395] = 12'hccc
rom[396] = 12'h777
rom[397] = 12'h777
rom[398] = 12'h777
rom[399] = 12'h777
rom[400] = 12'hfff
rom[401] = 12'hfff
rom[402] = 12'hfff
rom[403] = 12'hccc
rom[404] = 12'hccc
rom[405] = 12'hccc
rom[406] = 12'hccc
rom[407] = 12'hccc
rom[408] = 12'hccc
rom[409] = 12'hccc
rom[410] = 12'hccc
rom[411] = 12'hccc
rom[412] = 12'hccc
rom[413] = 12'hccc
rom[414] = 12'hccc
rom[415] = 12'hccc
rom[416] = 12'hccc
rom[417] = 12'hccc
rom[418] = 12'hccc
rom[419] = 12'hccc
rom[420] = 12'hccc
rom[421] = 12'h777
rom[422] = 12'h777
rom[423] = 12'h777
rom[424] = 12'h777
rom[425] = 12'hfff
rom[426] = 12'hfff
rom[427] = 12'hfff
rom[428] = 12'hccc
rom[429] = 12'hccc
rom[430] = 12'hccc
rom[431] = 12'hccc
rom[432] = 12'hccc
rom[433] = 12'hccc
rom[434] = 12'hccc
rom[435] = 12'hccc
rom[436] = 12'hccc
rom[437] = 12'hccc
rom[438] = 12'hccc
rom[439] = 12'hccc
rom[440] = 12'hbbb
rom[441] = 12'hccc
rom[442] = 12'hccc
rom[443] = 12'hccc
rom[444] = 12'hccc
rom[445] = 12'hccc
rom[446] = 12'h777
rom[447] = 12'h777
rom[448] = 12'h777
rom[449] = 12'h777
rom[450] = 12'hfff
rom[451] = 12'hfff
rom[452] = 12'hfff
rom[453] = 12'hccc
rom[454] = 12'hccc
rom[455] = 12'hccc
rom[456] = 12'hccc
rom[457] = 12'hccc
rom[458] = 12'hccc
rom[459] = 12'hccc
rom[460] = 12'hccc
rom[461] = 12'hccc
rom[462] = 12'hccc
rom[463] = 12'hccc
rom[464] = 12'hccc
rom[465] = 12'hbbb
rom[466] = 12'hccc
rom[467] = 12'hccc
rom[468] = 12'hccc
rom[469] = 12'hccc
rom[470] = 12'hccc
rom[471] = 12'h777
rom[472] = 12'h777
rom[473] = 12'h777
rom[474] = 12'h777
rom[475] = 12'hfff
rom[476] = 12'hfff
rom[477] = 12'hfff
rom[478] = 12'hccc
rom[479] = 12'hccc
rom[480] = 12'hccc
rom[481] = 12'hccc
rom[482] = 12'hccc
rom[483] = 12'hccc
rom[484] = 12'hccc
rom[485] = 12'hccc
rom[486] = 12'hccc
rom[487] = 12'hccc
rom[488] = 12'hccc
rom[489] = 12'hccc
rom[490] = 12'hccc
rom[491] = 12'hccc
rom[492] = 12'hccc
rom[493] = 12'hccc
rom[494] = 12'hccc
rom[495] = 12'hccc
rom[496] = 12'h777
rom[497] = 12'h777
rom[498] = 12'h777
rom[499] = 12'h777
rom[500] = 12'hfff
rom[501] = 12'hfff
rom[502] = 12'hfff
rom[503] = 12'hccc
rom[504] = 12'hccc
rom[505] = 12'hccc
rom[506] = 12'hccc
rom[507] = 12'hccc
rom[508] = 12'hccc
rom[509] = 12'hccc
rom[510] = 12'hccc
rom[511] = 12'hccc
rom[512] = 12'hccc
rom[513] = 12'hccc
rom[514] = 12'hccc
rom[515] = 12'hbbb
rom[516] = 12'hccc
rom[517] = 12'hccc
rom[518] = 12'hccc
rom[519] = 12'hccc
rom[520] = 12'hccc
rom[521] = 12'h777
rom[522] = 12'h777
rom[523] = 12'h777
rom[524] = 12'h777
rom[525] = 12'hfff
rom[526] = 12'hfff
rom[527] = 12'hfff
rom[528] = 12'h777
rom[529] = 12'h777
rom[530] = 12'h777
rom[531] = 12'h777
rom[532] = 12'h777
rom[533] = 12'h777
rom[534] = 12'h777
rom[535] = 12'h777
rom[536] = 12'h777
rom[537] = 12'h777
rom[538] = 12'h777
rom[539] = 12'h777
rom[540] = 12'h777
rom[541] = 12'h777
rom[542] = 12'h777
rom[543] = 12'h777
rom[544] = 12'h777
rom[545] = 12'h777
rom[546] = 12'h777
rom[547] = 12'h777
rom[548] = 12'h777
rom[549] = 12'h777
rom[550] = 12'hfff
rom[551] = 12'hfff
rom[552] = 12'h777
rom[553] = 12'h777
rom[554] = 12'h777
rom[555] = 12'h777
rom[556] = 12'h777
rom[557] = 12'h777
rom[558] = 12'h777
rom[559] = 12'h777
rom[560] = 12'h777
rom[561] = 12'h777
rom[562] = 12'h777
rom[563] = 12'h777
rom[564] = 12'h777
rom[565] = 12'h777
rom[566] = 12'h777
rom[567] = 12'h777
rom[568] = 12'h777
rom[569] = 12'h777
rom[570] = 12'h777
rom[571] = 12'h777
rom[572] = 12'h777
rom[573] = 12'h777
rom[574] = 12'h777
rom[575] = 12'hfff
rom[576] = 12'h777
rom[577] = 12'h777
rom[578] = 12'h777
rom[579] = 12'h777
rom[580] = 12'h777
rom[581] = 12'h777
rom[582] = 12'h777
rom[583] = 12'h777
rom[584] = 12'h777
rom[585] = 12'h777
rom[586] = 12'h777
rom[587] = 12'h777
rom[588] = 12'h777
rom[589] = 12'h777
rom[590] = 12'h777
rom[591] = 12'h777
rom[592] = 12'h777
rom[593] = 12'h777
rom[594] = 12'h777
rom[595] = 12'h888
rom[596] = 12'h777
rom[597] = 12'h777
rom[598] = 12'h777
rom[599] = 12'h777
rom[600] = 12'h777
rom[601] = 12'h777
rom[602] = 12'h777
rom[603] = 12'h777
rom[604] = 12'h777
rom[605] = 12'h777
rom[606] = 12'h777
rom[607] = 12'h777
rom[608] = 12'h777
rom[609] = 12'h777
rom[610] = 12'h777
rom[611] = 12'h777
rom[612] = 12'h777
rom[613] = 12'h777
rom[614] = 12'h777
rom[615] = 12'h777
rom[616] = 12'h777
rom[617] = 12'h777
rom[618] = 12'h777
rom[619] = 12'h777
rom[620] = 12'h777
rom[621] = 12'h777
rom[622] = 12'h777
rom[623] = 12'h777
rom[624] = 12'h777
  end

endmodule

module tile_flag_rom (                       //клетка с флагом
  input  wire    [13:0]     addr,
  output wire    [11:0]     word
);

  logic [11:0] rom [(25 * 25)];

  assign word = rom[addr];

  initial begin
rom[0] = 12'hfff
rom[1] = 12'hfff
rom[2] = 12'hfff
rom[3] = 12'hfff
rom[4] = 12'hfff
rom[5] = 12'hfff
rom[6] = 12'hfff
rom[7] = 12'hfff
rom[8] = 12'hfff
rom[9] = 12'hfff
rom[10] = 12'hfff
rom[11] = 12'hfff
rom[12] = 12'hfff
rom[13] = 12'hfff
rom[14] = 12'hfff
rom[15] = 12'hfff
rom[16] = 12'hfff
rom[17] = 12'hfff
rom[18] = 12'hfff
rom[19] = 12'hfff
rom[20] = 12'hfff
rom[21] = 12'hfff
rom[22] = 12'hfff
rom[23] = 12'hfff
rom[24] = 12'h777
rom[25] = 12'hfff
rom[26] = 12'hfff
rom[27] = 12'hfff
rom[28] = 12'hfff
rom[29] = 12'hfff
rom[30] = 12'hfff
rom[31] = 12'hfff
rom[32] = 12'hfff
rom[33] = 12'hfff
rom[34] = 12'hfff
rom[35] = 12'hfff
rom[36] = 12'hfff
rom[37] = 12'hfff
rom[38] = 12'hfff
rom[39] = 12'hfff
rom[40] = 12'hfff
rom[41] = 12'hfff
rom[42] = 12'hfff
rom[43] = 12'hfff
rom[44] = 12'hfff
rom[45] = 12'hfff
rom[46] = 12'hfff
rom[47] = 12'hfff
rom[48] = 12'h777
rom[49] = 12'h777
rom[50] = 12'hfff
rom[51] = 12'hfff
rom[52] = 12'hfff
rom[53] = 12'hfff
rom[54] = 12'hfff
rom[55] = 12'hfff
rom[56] = 12'hfff
rom[57] = 12'hfff
rom[58] = 12'hfff
rom[59] = 12'hfff
rom[60] = 12'hfff
rom[61] = 12'hfff
rom[62] = 12'hfff
rom[63] = 12'hfff
rom[64] = 12'hfff
rom[65] = 12'hfff
rom[66] = 12'hfff
rom[67] = 12'hfff
rom[68] = 12'hfff
rom[69] = 12'hfff
rom[70] = 12'hfff
rom[71] = 12'hfff
rom[72] = 12'h777
rom[73] = 12'h777
rom[74] = 12'h777
rom[75] = 12'hfff
rom[76] = 12'hfff
rom[77] = 12'hfff
rom[78] = 12'hccc
rom[79] = 12'hccc
rom[80] = 12'hccc
rom[81] = 12'hccc
rom[82] = 12'hccc
rom[83] = 12'hccc
rom[84] = 12'hccc
rom[85] = 12'hccc
rom[86] = 12'hccc
rom[87] = 12'hccc
rom[88] = 12'hccc
rom[89] = 12'hccc
rom[90] = 12'hccc
rom[91] = 12'hccc
rom[92] = 12'hccc
rom[93] = 12'hccc
rom[94] = 12'hccc
rom[95] = 12'hccc
rom[96] = 12'h777
rom[97] = 12'h777
rom[98] = 12'h777
rom[99] = 12'h777
rom[100] = 12'hfff
rom[101] = 12'hfff
rom[102] = 12'hfff
rom[103] = 12'hccc
rom[104] = 12'hccc
rom[105] = 12'hccc
rom[106] = 12'hccc
rom[107] = 12'hccc
rom[108] = 12'hccc
rom[109] = 12'hccc
rom[110] = 12'hccc
rom[111] = 12'hccc
rom[112] = 12'hccc
rom[113] = 12'hccc
rom[114] = 12'hccc
rom[115] = 12'hccc
rom[116] = 12'hccc
rom[117] = 12'hccc
rom[118] = 12'hccc
rom[119] = 12'hccc
rom[120] = 12'hccc
rom[121] = 12'h777
rom[122] = 12'h777
rom[123] = 12'h777
rom[124] = 12'h777
rom[125] = 12'hfff
rom[126] = 12'hfff
rom[127] = 12'hfff
rom[128] = 12'hccc
rom[129] = 12'hccc
rom[130] = 12'hccc
rom[131] = 12'hccc
rom[132] = 12'hccc
rom[133] = 12'hccc
rom[134] = 12'hccc
rom[135] = 12'hccc
rom[136] = 12'hccc
rom[137] = 12'hccc
rom[138] = 12'hccc
rom[139] = 12'hccc
rom[140] = 12'hccc
rom[141] = 12'hccc
rom[142] = 12'hccc
rom[143] = 12'hccc
rom[144] = 12'hccc
rom[145] = 12'hccc
rom[146] = 12'h777
rom[147] = 12'h777
rom[148] = 12'h777
rom[149] = 12'h777
rom[150] = 12'hfff
rom[151] = 12'hfff
rom[152] = 12'hfff
rom[153] = 12'hccc
rom[154] = 12'hccc
rom[155] = 12'hccc
rom[156] = 12'hccc
rom[157] = 12'hccc
rom[158] = 12'hccc
rom[159] = 12'hccc
rom[160] = 12'hccc
rom[161] = 12'hccc
rom[162] = 12'hccc
rom[163] = 12'hccc
rom[164] = 12'hccc
rom[165] = 12'hccc
rom[166] = 12'hccc
rom[167] = 12'hccc
rom[168] = 12'hccc
rom[169] = 12'hccc
rom[170] = 12'hccc
rom[171] = 12'h777
rom[172] = 12'h777
rom[173] = 12'h777
rom[174] = 12'h777
rom[175] = 12'hfff
rom[176] = 12'hfff
rom[177] = 12'hfff
rom[178] = 12'hccc
rom[179] = 12'hccc
rom[180] = 12'hccc
rom[181] = 12'hccc
rom[182] = 12'hccc
rom[183] = 12'hccc
rom[184] = 12'hccc
rom[185] = 12'hccc
rom[186] = 12'h00f
rom[187] = 12'h00f
rom[188] = 12'hccc
rom[189] = 12'hccc
rom[190] = 12'hccc
rom[191] = 12'hccc
rom[192] = 12'hccc
rom[193] = 12'hccc
rom[194] = 12'hccc
rom[195] = 12'hccc
rom[196] = 12'h777
rom[197] = 12'h777
rom[198] = 12'h777
rom[199] = 12'h777
rom[200] = 12'hfff
rom[201] = 12'hfff
rom[202] = 12'hfff
rom[203] = 12'hccc
rom[204] = 12'hccc
rom[205] = 12'hccc
rom[206] = 12'hccc
rom[207] = 12'hccc
rom[208] = 12'hccc
rom[209] = 12'h00f
rom[210] = 12'h00f
rom[211] = 12'h00f
rom[212] = 12'h00f
rom[213] = 12'hccc
rom[214] = 12'hccc
rom[215] = 12'hccc
rom[216] = 12'hccc
rom[217] = 12'hccc
rom[218] = 12'hccc
rom[219] = 12'hccc
rom[220] = 12'hccc
rom[221] = 12'h777
rom[222] = 12'h777
rom[223] = 12'h777
rom[224] = 12'h777
rom[225] = 12'hfff
rom[226] = 12'hfff
rom[227] = 12'hfff
rom[228] = 12'hccc
rom[229] = 12'hccc
rom[230] = 12'hccc
rom[231] = 12'hccc
rom[232] = 12'hccc
rom[233] = 12'h00f
rom[234] = 12'h00f
rom[235] = 12'h00f
rom[236] = 12'h00f
rom[237] = 12'h00f
rom[238] = 12'hccc
rom[239] = 12'hccc
rom[240] = 12'hccc
rom[241] = 12'hccc
rom[242] = 12'hccc
rom[243] = 12'hccc
rom[244] = 12'hccc
rom[245] = 12'hccc
rom[246] = 12'h777
rom[247] = 12'h777
rom[248] = 12'h777
rom[249] = 12'h777
rom[250] = 12'hfff
rom[251] = 12'hfff
rom[252] = 12'hfff
rom[253] = 12'hccc
rom[254] = 12'hccc
rom[255] = 12'hccc
rom[256] = 12'hccc
rom[257] = 12'hccc
rom[258] = 12'hccc
rom[259] = 12'h00f
rom[260] = 12'h00f
rom[261] = 12'h00f
rom[262] = 12'h00f
rom[263] = 12'hccc
rom[264] = 12'hccc
rom[265] = 12'hccc
rom[266] = 12'hccc
rom[267] = 12'hccc
rom[268] = 12'hccc
rom[269] = 12'hccc
rom[270] = 12'hccc
rom[271] = 12'h777
rom[272] = 12'h777
rom[273] = 12'h777
rom[274] = 12'h777
rom[275] = 12'hfff
rom[276] = 12'hfff
rom[277] = 12'hfff
rom[278] = 12'hccc
rom[279] = 12'hccc
rom[280] = 12'hccc
rom[281] = 12'hccc
rom[282] = 12'hccc
rom[283] = 12'hccc
rom[284] = 12'hccc
rom[285] = 12'hccc
rom[286] = 12'h00f
rom[287] = 12'h00f
rom[288] = 12'hccc
rom[289] = 12'hccc
rom[290] = 12'hccc
rom[291] = 12'hccc
rom[292] = 12'hccc
rom[293] = 12'hccc
rom[294] = 12'hccc
rom[295] = 12'hccc
rom[296] = 12'h777
rom[297] = 12'h777
rom[298] = 12'h777
rom[299] = 12'h777
rom[300] = 12'hfff
rom[301] = 12'hfff
rom[302] = 12'hfff
rom[303] = 12'hccc
rom[304] = 12'hccc
rom[305] = 12'hccc
rom[306] = 12'hccc
rom[307] = 12'hccc
rom[308] = 12'hccc
rom[309] = 12'hccc
rom[310] = 12'hccc
rom[311] = 12'hccc
rom[312] = 12'h000
rom[313] = 12'hccc
rom[314] = 12'hccc
rom[315] = 12'hccc
rom[316] = 12'hccc
rom[317] = 12'hccc
rom[318] = 12'hccc
rom[319] = 12'hccc
rom[320] = 12'hccc
rom[321] = 12'h777
rom[322] = 12'h777
rom[323] = 12'h777
rom[324] = 12'h777
rom[325] = 12'hfff
rom[326] = 12'hfff
rom[327] = 12'hfff
rom[328] = 12'hccc
rom[329] = 12'hccc
rom[330] = 12'hccc
rom[331] = 12'hccc
rom[332] = 12'hccc
rom[333] = 12'hccc
rom[334] = 12'hccc
rom[335] = 12'hccc
rom[336] = 12'hccc
rom[337] = 12'h000
rom[338] = 12'hccc
rom[339] = 12'hccc
rom[340] = 12'hccc
rom[341] = 12'hccc
rom[342] = 12'hccc
rom[343] = 12'hccc
rom[344] = 12'hccc
rom[345] = 12'hccc
rom[346] = 12'h777
rom[347] = 12'h777
rom[348] = 12'h777
rom[349] = 12'h777
rom[350] = 12'hfff
rom[351] = 12'hfff
rom[352] = 12'hfff
rom[353] = 12'hccc
rom[354] = 12'hccc
rom[355] = 12'hccc
rom[356] = 12'hccc
rom[357] = 12'hccc
rom[358] = 12'hccc
rom[359] = 12'hccc
rom[360] = 12'h000
rom[361] = 12'h000
rom[362] = 12'h000
rom[363] = 12'h000
rom[364] = 12'hccc
rom[365] = 12'hccc
rom[366] = 12'hccc
rom[367] = 12'hccc
rom[368] = 12'hccc
rom[369] = 12'hccc
rom[370] = 12'hccc
rom[371] = 12'h777
rom[372] = 12'h777
rom[373] = 12'h777
rom[374] = 12'h777
rom[375] = 12'hfff
rom[376] = 12'hfff
rom[377] = 12'hfff
rom[378] = 12'hccc
rom[379] = 12'hccc
rom[380] = 12'hccc
rom[381] = 12'hccc
rom[382] = 12'hccc
rom[383] = 12'h000
rom[384] = 12'h000
rom[385] = 12'h000
rom[386] = 12'h000
rom[387] = 12'h000
rom[388] = 12'h000
rom[389] = 12'h000
rom[390] = 12'h000
rom[391] = 12'hccc
rom[392] = 12'hccc
rom[393] = 12'hccc
rom[394] = 12'hccc
rom[395] = 12'hccc
rom[396] = 12'h777
rom[397] = 12'h777
rom[398] = 12'h777
rom[399] = 12'h777
rom[400] = 12'hfff
rom[401] = 12'hfff
rom[402] = 12'hfff
rom[403] = 12'hccc
rom[404] = 12'hccc
rom[405] = 12'hccc
rom[406] = 12'hccc
rom[407] = 12'hccc
rom[408] = 12'h000
rom[409] = 12'h000
rom[410] = 12'h000
rom[411] = 12'h000
rom[412] = 12'h000
rom[413] = 12'h000
rom[414] = 12'h000
rom[415] = 12'h000
rom[416] = 12'hccc
rom[417] = 12'hccc
rom[418] = 12'hccc
rom[419] = 12'hccc
rom[420] = 12'hccc
rom[421] = 12'h777
rom[422] = 12'h777
rom[423] = 12'h777
rom[424] = 12'h777
rom[425] = 12'hfff
rom[426] = 12'hfff
rom[427] = 12'hfff
rom[428] = 12'hccc
rom[429] = 12'hccc
rom[430] = 12'hccc
rom[431] = 12'hccc
rom[432] = 12'hccc
rom[433] = 12'hccc
rom[434] = 12'hccc
rom[435] = 12'hccc
rom[436] = 12'hccc
rom[437] = 12'hccc
rom[438] = 12'hccc
rom[439] = 12'hccc
rom[440] = 12'hbbb
rom[441] = 12'hccc
rom[442] = 12'hccc
rom[443] = 12'hccc
rom[444] = 12'hccc
rom[445] = 12'hccc
rom[446] = 12'h777
rom[447] = 12'h777
rom[448] = 12'h777
rom[449] = 12'h777
rom[450] = 12'hfff
rom[451] = 12'hfff
rom[452] = 12'hfff
rom[453] = 12'hccc
rom[454] = 12'hccc
rom[455] = 12'hccc
rom[456] = 12'hccc
rom[457] = 12'hccc
rom[458] = 12'hccc
rom[459] = 12'hccc
rom[460] = 12'hccc
rom[461] = 12'hccc
rom[462] = 12'hccc
rom[463] = 12'hccc
rom[464] = 12'hccc
rom[465] = 12'hbbb
rom[466] = 12'hccc
rom[467] = 12'hccc
rom[468] = 12'hccc
rom[469] = 12'hccc
rom[470] = 12'hccc
rom[471] = 12'h777
rom[472] = 12'h777
rom[473] = 12'h777
rom[474] = 12'h777
rom[475] = 12'hfff
rom[476] = 12'hfff
rom[477] = 12'hfff
rom[478] = 12'hccc
rom[479] = 12'hccc
rom[480] = 12'hccc
rom[481] = 12'hccc
rom[482] = 12'hccc
rom[483] = 12'hccc
rom[484] = 12'hccc
rom[485] = 12'hccc
rom[486] = 12'hccc
rom[487] = 12'hccc
rom[488] = 12'hccc
rom[489] = 12'hccc
rom[490] = 12'hccc
rom[491] = 12'hccc
rom[492] = 12'hccc
rom[493] = 12'hccc
rom[494] = 12'hccc
rom[495] = 12'hccc
rom[496] = 12'h777
rom[497] = 12'h777
rom[498] = 12'h777
rom[499] = 12'h777
rom[500] = 12'hfff
rom[501] = 12'hfff
rom[502] = 12'hfff
rom[503] = 12'hccc
rom[504] = 12'hccc
rom[505] = 12'hccc
rom[506] = 12'hccc
rom[507] = 12'hccc
rom[508] = 12'hccc
rom[509] = 12'hccc
rom[510] = 12'hccc
rom[511] = 12'hccc
rom[512] = 12'hccc
rom[513] = 12'hccc
rom[514] = 12'hccc
rom[515] = 12'hbbb
rom[516] = 12'hccc
rom[517] = 12'hccc
rom[518] = 12'hccc
rom[519] = 12'hccc
rom[520] = 12'hccc
rom[521] = 12'h777
rom[522] = 12'h777
rom[523] = 12'h777
rom[524] = 12'h777
rom[525] = 12'hfff
rom[526] = 12'hfff
rom[527] = 12'hfff
rom[528] = 12'h777
rom[529] = 12'h777
rom[530] = 12'h777
rom[531] = 12'h777
rom[532] = 12'h777
rom[533] = 12'h777
rom[534] = 12'h777
rom[535] = 12'h777
rom[536] = 12'h777
rom[537] = 12'h777
rom[538] = 12'h777
rom[539] = 12'h777
rom[540] = 12'h777
rom[541] = 12'h777
rom[542] = 12'h777
rom[543] = 12'h777
rom[544] = 12'h777
rom[545] = 12'h777
rom[546] = 12'h777
rom[547] = 12'h777
rom[548] = 12'h777
rom[549] = 12'h777
rom[550] = 12'hfff
rom[551] = 12'hfff
rom[552] = 12'h777
rom[553] = 12'h777
rom[554] = 12'h777
rom[555] = 12'h777
rom[556] = 12'h777
rom[557] = 12'h777
rom[558] = 12'h777
rom[559] = 12'h777
rom[560] = 12'h777
rom[561] = 12'h777
rom[562] = 12'h777
rom[563] = 12'h777
rom[564] = 12'h777
rom[565] = 12'h777
rom[566] = 12'h777
rom[567] = 12'h777
rom[568] = 12'h777
rom[569] = 12'h777
rom[570] = 12'h777
rom[571] = 12'h777
rom[572] = 12'h777
rom[573] = 12'h777
rom[574] = 12'h777
rom[575] = 12'hfff
rom[576] = 12'h777
rom[577] = 12'h777
rom[578] = 12'h777
rom[579] = 12'h777
rom[580] = 12'h777
rom[581] = 12'h777
rom[582] = 12'h777
rom[583] = 12'h777
rom[584] = 12'h777
rom[585] = 12'h777
rom[586] = 12'h777
rom[587] = 12'h777
rom[588] = 12'h777
rom[589] = 12'h777
rom[590] = 12'h777
rom[591] = 12'h777
rom[592] = 12'h777
rom[593] = 12'h777
rom[594] = 12'h777
rom[595] = 12'h888
rom[596] = 12'h777
rom[597] = 12'h777
rom[598] = 12'h777
rom[599] = 12'h777
rom[600] = 12'h777
rom[601] = 12'h777
rom[602] = 12'h777
rom[603] = 12'h777
rom[604] = 12'h777
rom[605] = 12'h777
rom[606] = 12'h777
rom[607] = 12'h777
rom[608] = 12'h777
rom[609] = 12'h777
rom[610] = 12'h777
rom[611] = 12'h777
rom[612] = 12'h777
rom[613] = 12'h777
rom[614] = 12'h777
rom[615] = 12'h777
rom[616] = 12'h777
rom[617] = 12'h777
rom[618] = 12'h777
rom[619] = 12'h777
rom[620] = 12'h777
rom[621] = 12'h777
rom[622] = 12'h777
rom[623] = 12'h777
rom[624] = 12'h777
  end
endmodule

module tile_one_rom (                       //клетка с единицей
  input  wire    [13:0]     addr,
  output wire    [11:0]     word
);

  logic [11:0] rom [(25 * 25)];

  assign word = rom[addr];

  initial begin
rom[0] = 12'h777;
rom[1] = 12'h777;
rom[2] = 12'h777;
rom[3] = 12'h777;
rom[4] = 12'h777;
rom[5] = 12'h777;
rom[6] = 12'h777;
rom[7] = 12'h777;
rom[8] = 12'h777;
rom[9] = 12'h777;
rom[10] = 12'h777;
rom[11] = 12'h777;
rom[12] = 12'h777;
rom[13] = 12'h777;
rom[14] = 12'h777;
rom[15] = 12'h777;
rom[16] = 12'h777;
rom[17] = 12'h777;
rom[18] = 12'h777;
rom[19] = 12'h777;
rom[20] = 12'h777;
rom[21] = 12'h777;
rom[22] = 12'h777;
rom[23] = 12'h777;
rom[24] = 12'h777;
rom[25] = 12'h777;
rom[26] = 12'hccc;
rom[27] = 12'hccc;
rom[28] = 12'hccc;
rom[29] = 12'hccc;
rom[30] = 12'hccc;
rom[31] = 12'hccc;
rom[32] = 12'hccc;
rom[33] = 12'hccc;
rom[34] = 12'hccc;
rom[35] = 12'hccc;
rom[36] = 12'hccc;
rom[37] = 12'hccc;
rom[38] = 12'hccc;
rom[39] = 12'hccc;
rom[40] = 12'hccc;
rom[41] = 12'hccc;
rom[42] = 12'hccc;
rom[43] = 12'hccc;
rom[44] = 12'hccc;
rom[45] = 12'hccc;
rom[46] = 12'hccc;
rom[47] = 12'hccc;
rom[48] = 12'hccc;
rom[49] = 12'h777;
rom[50] = 12'h777;
rom[51] = 12'hccc;
rom[52] = 12'hccc;
rom[53] = 12'hccc;
rom[54] = 12'hccc;
rom[55] = 12'hccc;
rom[56] = 12'hccc;
rom[57] = 12'hccc;
rom[58] = 12'hccc;
rom[59] = 12'hccc;
rom[60] = 12'hccc;
rom[61] = 12'hccc;
rom[62] = 12'hccc;
rom[63] = 12'hccc;
rom[64] = 12'hccc;
rom[65] = 12'hccc;
rom[66] = 12'hccc;
rom[67] = 12'hccc;
rom[68] = 12'hccc;
rom[69] = 12'hccc;
rom[70] = 12'hccc;
rom[71] = 12'hccc;
rom[72] = 12'hccc;
rom[73] = 12'hccc;
rom[74] = 12'h777;
rom[75] = 12'h777;
rom[76] = 12'hccc;
rom[77] = 12'hccc;
rom[78] = 12'hccc;
rom[79] = 12'hccc;
rom[80] = 12'hccc;
rom[81] = 12'hccc;
rom[82] = 12'hccc;
rom[83] = 12'hccc;
rom[84] = 12'hccc;
rom[85] = 12'hccc;
rom[86] = 12'hccc;
rom[87] = 12'hccc;
rom[88] = 12'hccc;
rom[89] = 12'hccc;
rom[90] = 12'hccc;
rom[91] = 12'hccc;
rom[92] = 12'hccc;
rom[93] = 12'hccc;
rom[94] = 12'hccc;
rom[95] = 12'hccc;
rom[96] = 12'hccc;
rom[97] = 12'hccc;
rom[98] = 12'hccc;
rom[99] = 12'h777;
rom[100] = 12'h777;
rom[101] = 12'hccc;
rom[102] = 12'hccc;
rom[103] = 12'hccc;
rom[104] = 12'hccc;
rom[105] = 12'hccc;
rom[106] = 12'hccc;
rom[107] = 12'hccc;
rom[108] = 12'hccc;
rom[109] = 12'hccc;
rom[110] = 12'hccc;
rom[111] = 12'hccc;
rom[112] = 12'hccc;
rom[113] = 12'hccc;
rom[114] = 12'hccc;
rom[115] = 12'hccc;
rom[116] = 12'hccc;
rom[117] = 12'hccc;
rom[118] = 12'hccc;
rom[119] = 12'hccc;
rom[120] = 12'hccc;
rom[121] = 12'hccc;
rom[122] = 12'hccc;
rom[123] = 12'hccc;
rom[124] = 12'h777;
rom[125] = 12'h777;
rom[126] = 12'hccc;
rom[127] = 12'hccc;
rom[128] = 12'hccc;
rom[129] = 12'hccc;
rom[130] = 12'hccc;
rom[131] = 12'hccc;
rom[132] = 12'hccc;
rom[133] = 12'hccc;
rom[134] = 12'hccc;
rom[135] = 12'hccc;
rom[136] = 12'hccc;
rom[137] = 12'hccc;
rom[138] = 12'hccc;
rom[139] = 12'hccc;
rom[140] = 12'hccc;
rom[141] = 12'hccc;
rom[142] = 12'hccc;
rom[143] = 12'hccc;
rom[144] = 12'hccc;
rom[145] = 12'hccc;
rom[146] = 12'hccc;
rom[147] = 12'hccc;
rom[148] = 12'hccc;
rom[149] = 12'h777;
rom[150] = 12'h777;
rom[151] = 12'hccc;
rom[152] = 12'hccc;
rom[153] = 12'hccc;
rom[154] = 12'hccc;
rom[155] = 12'hccc;
rom[156] = 12'hccc;
rom[157] = 12'hccc;
rom[158] = 12'hccc;
rom[159] = 12'hccc;
rom[160] = 12'hccc;
rom[161] = 12'hccc;
rom[162] = 12'hccc;
rom[163] = 12'hccc;
rom[164] = 12'hccc;
rom[165] = 12'hccc;
rom[166] = 12'hccc;
rom[167] = 12'hccc;
rom[168] = 12'hccc;
rom[169] = 12'hccc;
rom[170] = 12'hccc;
rom[171] = 12'hccc;
rom[172] = 12'hccc;
rom[173] = 12'hccc;
rom[174] = 12'h777;
rom[175] = 12'h777;
rom[176] = 12'hccc;
rom[177] = 12'hccc;
rom[178] = 12'hccc;
rom[179] = 12'hccc;
rom[180] = 12'hccc;
rom[181] = 12'hccc;
rom[182] = 12'hccc;
rom[183] = 12'hccc;
rom[184] = 12'hccc;
rom[185] = 12'hccc;
rom[186] = 12'hccc;
rom[187] = 12'hf00;
rom[188] = 12'hf00;
rom[189] = 12'hccc;
rom[190] = 12'hccc;
rom[191] = 12'hccc;
rom[192] = 12'hccc;
rom[193] = 12'hccc;
rom[194] = 12'hccc;
rom[195] = 12'hccc;
rom[196] = 12'hccc;
rom[197] = 12'hccc;
rom[198] = 12'hccc;
rom[199] = 12'h777;
rom[200] = 12'h777;
rom[201] = 12'hccc;
rom[202] = 12'hccc;
rom[203] = 12'hccc;
rom[204] = 12'hccc;
rom[205] = 12'hccc;
rom[206] = 12'hccc;
rom[207] = 12'hccc;
rom[208] = 12'hccc;
rom[209] = 12'hccc;
rom[210] = 12'hccc;
rom[211] = 12'hf00;
rom[212] = 12'hf00;
rom[213] = 12'hf00;
rom[214] = 12'hccc;
rom[215] = 12'hccc;
rom[216] = 12'hccc;
rom[217] = 12'hccc;
rom[218] = 12'hccc;
rom[219] = 12'hccc;
rom[220] = 12'hccc;
rom[221] = 12'hccc;
rom[222] = 12'hccc;
rom[223] = 12'hccc;
rom[224] = 12'h777;
rom[225] = 12'h777;
rom[226] = 12'hccc;
rom[227] = 12'hccc;
rom[228] = 12'hccc;
rom[229] = 12'hccc;
rom[230] = 12'hccc;
rom[231] = 12'hccc;
rom[232] = 12'hccc;
rom[233] = 12'hccc;
rom[234] = 12'hccc;
rom[235] = 12'hf00;
rom[236] = 12'hf00;
rom[237] = 12'hf00;
rom[238] = 12'hf00;
rom[239] = 12'hccc;
rom[240] = 12'hccc;
rom[241] = 12'hccc;
rom[242] = 12'hccc;
rom[243] = 12'hccc;
rom[244] = 12'hccc;
rom[245] = 12'hccc;
rom[246] = 12'hccc;
rom[247] = 12'hccc;
rom[248] = 12'hccc;
rom[249] = 12'h777;
rom[250] = 12'h777;
rom[251] = 12'hccc;
rom[252] = 12'hccc;
rom[253] = 12'hccc;
rom[254] = 12'hccc;
rom[255] = 12'hccc;
rom[256] = 12'hccc;
rom[257] = 12'hccc;
rom[258] = 12'hccc;
rom[259] = 12'hf00;
rom[260] = 12'hf00;
rom[261] = 12'hf00;
rom[262] = 12'hf00;
rom[263] = 12'hf00;
rom[264] = 12'hccc;
rom[265] = 12'hccc;
rom[266] = 12'hccc;
rom[267] = 12'hccc;
rom[268] = 12'hccc;
rom[269] = 12'hccc;
rom[270] = 12'hccc;
rom[271] = 12'hccc;
rom[272] = 12'hccc;
rom[273] = 12'hccc;
rom[274] = 12'h777;
rom[275] = 12'h777;
rom[276] = 12'hccc;
rom[277] = 12'hccc;
rom[278] = 12'hccc;
rom[279] = 12'hccc;
rom[280] = 12'hccc;
rom[281] = 12'hccc;
rom[282] = 12'hccc;
rom[283] = 12'hccc;
rom[284] = 12'hccc;
rom[285] = 12'hccc;
rom[286] = 12'hf00;
rom[287] = 12'hf00;
rom[288] = 12'hf00;
rom[289] = 12'hccc;
rom[290] = 12'hccc;
rom[291] = 12'hccc;
rom[292] = 12'hccc;
rom[293] = 12'hccc;
rom[294] = 12'hccc;
rom[295] = 12'hccc;
rom[296] = 12'hccc;
rom[297] = 12'hccc;
rom[298] = 12'hccc;
rom[299] = 12'h777;
rom[300] = 12'h777;
rom[301] = 12'hccc;
rom[302] = 12'hccc;
rom[303] = 12'hccc;
rom[304] = 12'hccc;
rom[305] = 12'hccc;
rom[306] = 12'hccc;
rom[307] = 12'hccc;
rom[308] = 12'hccc;
rom[309] = 12'hccc;
rom[310] = 12'hccc;
rom[311] = 12'hf00;
rom[312] = 12'hf00;
rom[313] = 12'hf00;
rom[314] = 12'hccc;
rom[315] = 12'hccc;
rom[316] = 12'hccc;
rom[317] = 12'hccc;
rom[318] = 12'hccc;
rom[319] = 12'hccc;
rom[320] = 12'hccc;
rom[321] = 12'hccc;
rom[322] = 12'hccc;
rom[323] = 12'hccc;
rom[324] = 12'h777;
rom[325] = 12'h777;
rom[326] = 12'hccc;
rom[327] = 12'hccc;
rom[328] = 12'hccc;
rom[329] = 12'hccc;
rom[330] = 12'hccc;
rom[331] = 12'hccc;
rom[332] = 12'hccc;
rom[333] = 12'hccc;
rom[334] = 12'hccc;
rom[335] = 12'hccc;
rom[336] = 12'hf00;
rom[337] = 12'hf00;
rom[338] = 12'hf00;
rom[339] = 12'hccc;
rom[340] = 12'hccc;
rom[341] = 12'hccc;
rom[342] = 12'hccc;
rom[343] = 12'hccc;
rom[344] = 12'hccc;
rom[345] = 12'hccc;
rom[346] = 12'hccc;
rom[347] = 12'hccc;
rom[348] = 12'hccc;
rom[349] = 12'h777;
rom[350] = 12'h777;
rom[351] = 12'hccc;
rom[352] = 12'hccc;
rom[353] = 12'hccc;
rom[354] = 12'hccc;
rom[355] = 12'hccc;
rom[356] = 12'hccc;
rom[357] = 12'hccc;
rom[358] = 12'hccc;
rom[359] = 12'hccc;
rom[360] = 12'hccc;
rom[361] = 12'hf00;
rom[362] = 12'hf00;
rom[363] = 12'hf00;
rom[364] = 12'hccc;
rom[365] = 12'hccc;
rom[366] = 12'hccc;
rom[367] = 12'hccc;
rom[368] = 12'hccc;
rom[369] = 12'hccc;
rom[370] = 12'hccc;
rom[371] = 12'hccc;
rom[372] = 12'hccc;
rom[373] = 12'hccc;
rom[374] = 12'h777;
rom[375] = 12'h777;
rom[376] = 12'hccc;
rom[377] = 12'hccc;
rom[378] = 12'hccc;
rom[379] = 12'hccc;
rom[380] = 12'hccc;
rom[381] = 12'hccc;
rom[382] = 12'hccc;
rom[383] = 12'hccc;
rom[384] = 12'hf00;
rom[385] = 12'hf00;
rom[386] = 12'hf00;
rom[387] = 12'hf00;
rom[388] = 12'hf00;
rom[389] = 12'hf00;
rom[390] = 12'hf00;
rom[391] = 12'hccc;
rom[392] = 12'hccc;
rom[393] = 12'hccc;
rom[394] = 12'hccc;
rom[395] = 12'hccc;
rom[396] = 12'hccc;
rom[397] = 12'hccc;
rom[398] = 12'hccc;
rom[399] = 12'h777;
rom[400] = 12'h777;
rom[401] = 12'hccc;
rom[402] = 12'hccc;
rom[403] = 12'hccc;
rom[404] = 12'hccc;
rom[405] = 12'hccc;
rom[406] = 12'hccc;
rom[407] = 12'hccc;
rom[408] = 12'hccc;
rom[409] = 12'hf00;
rom[410] = 12'hf00;
rom[411] = 12'hf00;
rom[412] = 12'hf00;
rom[413] = 12'hf00;
rom[414] = 12'hf00;
rom[415] = 12'hf00;
rom[416] = 12'hccc;
rom[417] = 12'hccc;
rom[418] = 12'hccc;
rom[419] = 12'hccc;
rom[420] = 12'hccc;
rom[421] = 12'hccc;
rom[422] = 12'hccc;
rom[423] = 12'hccc;
rom[424] = 12'h777;
rom[425] = 12'h777;
rom[426] = 12'hccc;
rom[427] = 12'hccc;
rom[428] = 12'hccc;
rom[429] = 12'hccc;
rom[430] = 12'hccc;
rom[431] = 12'hccc;
rom[432] = 12'hccc;
rom[433] = 12'hccc;
rom[434] = 12'hccc;
rom[435] = 12'hccc;
rom[436] = 12'hccc;
rom[437] = 12'hccc;
rom[438] = 12'hccc;
rom[439] = 12'hccc;
rom[440] = 12'hbbb;
rom[441] = 12'hccc;
rom[442] = 12'hccc;
rom[443] = 12'hccc;
rom[444] = 12'hccc;
rom[445] = 12'hccc;
rom[446] = 12'hccc;
rom[447] = 12'hccc;
rom[448] = 12'hccc;
rom[449] = 12'h777;
rom[450] = 12'h777;
rom[451] = 12'hccc;
rom[452] = 12'hccc;
rom[453] = 12'hccc;
rom[454] = 12'hccc;
rom[455] = 12'hccc;
rom[456] = 12'hccc;
rom[457] = 12'hccc;
rom[458] = 12'hccc;
rom[459] = 12'hccc;
rom[460] = 12'hccc;
rom[461] = 12'hccc;
rom[462] = 12'hccc;
rom[463] = 12'hccc;
rom[464] = 12'hccc;
rom[465] = 12'hbbb;
rom[466] = 12'hccc;
rom[467] = 12'hccc;
rom[468] = 12'hccc;
rom[469] = 12'hccc;
rom[470] = 12'hccc;
rom[471] = 12'hccc;
rom[472] = 12'hccc;
rom[473] = 12'hccc;
rom[474] = 12'h777;
rom[475] = 12'h777;
rom[476] = 12'hccc;
rom[477] = 12'hccc;
rom[478] = 12'hccc;
rom[479] = 12'hccc;
rom[480] = 12'hccc;
rom[481] = 12'hccc;
rom[482] = 12'hccc;
rom[483] = 12'hccc;
rom[484] = 12'hccc;
rom[485] = 12'hccc;
rom[486] = 12'hccc;
rom[487] = 12'hccc;
rom[488] = 12'hccc;
rom[489] = 12'hccc;
rom[490] = 12'hccc;
rom[491] = 12'hccc;
rom[492] = 12'hccc;
rom[493] = 12'hccc;
rom[494] = 12'hccc;
rom[495] = 12'hccc;
rom[496] = 12'hccc;
rom[497] = 12'hccc;
rom[498] = 12'hccc;
rom[499] = 12'h777;
rom[500] = 12'h777;
rom[501] = 12'hccc;
rom[502] = 12'hccc;
rom[503] = 12'hccc;
rom[504] = 12'hccc;
rom[505] = 12'hccc;
rom[506] = 12'hccc;
rom[507] = 12'hccc;
rom[508] = 12'hccc;
rom[509] = 12'hccc;
rom[510] = 12'hccc;
rom[511] = 12'hccc;
rom[512] = 12'hccc;
rom[513] = 12'hccc;
rom[514] = 12'hccc;
rom[515] = 12'hccc;
rom[516] = 12'hccc;
rom[517] = 12'hccc;
rom[518] = 12'hccc;
rom[519] = 12'hccc;
rom[520] = 12'hccc;
rom[521] = 12'hccc;
rom[522] = 12'hccc;
rom[523] = 12'hccc;
rom[524] = 12'h777;
rom[525] = 12'h777;
rom[526] = 12'hccc;
rom[527] = 12'hccc;
rom[528] = 12'hccc;
rom[529] = 12'hccc;
rom[530] = 12'hccc;
rom[531] = 12'hccc;
rom[532] = 12'hccc;
rom[533] = 12'hccc;
rom[534] = 12'hccc;
rom[535] = 12'hccc;
rom[536] = 12'hccc;
rom[537] = 12'hccc;
rom[538] = 12'hccc;
rom[539] = 12'hccc;
rom[540] = 12'hccc;
rom[541] = 12'hccc;
rom[542] = 12'hccc;
rom[543] = 12'hccc;
rom[544] = 12'hccc;
rom[545] = 12'hccc;
rom[546] = 12'hccc;
rom[547] = 12'hccc;
rom[548] = 12'hccc;
rom[549] = 12'h777;
rom[550] = 12'h777;
rom[551] = 12'hccc;
rom[552] = 12'hccc;
rom[553] = 12'hccc;
rom[554] = 12'hccc;
rom[555] = 12'hccc;
rom[556] = 12'hccc;
rom[557] = 12'hccc;
rom[558] = 12'hccc;
rom[559] = 12'hccc;
rom[560] = 12'hccc;
rom[561] = 12'hccc;
rom[562] = 12'hccc;
rom[563] = 12'hccc;
rom[564] = 12'hccc;
rom[565] = 12'hccc;
rom[566] = 12'hccc;
rom[567] = 12'hccc;
rom[568] = 12'hccc;
rom[569] = 12'hccc;
rom[570] = 12'hccc;
rom[571] = 12'hccc;
rom[572] = 12'hccc;
rom[573] = 12'hccc;
rom[574] = 12'h777;
rom[575] = 12'h777;
rom[576] = 12'hccc;
rom[577] = 12'hccc;
rom[578] = 12'hccc;
rom[579] = 12'hccc;
rom[580] = 12'hccc;
rom[581] = 12'hccc;
rom[582] = 12'hccc;
rom[583] = 12'hccc;
rom[584] = 12'hccc;
rom[585] = 12'hccc;
rom[586] = 12'hccc;
rom[587] = 12'hccc;
rom[588] = 12'hccc;
rom[589] = 12'hccc;
rom[590] = 12'hccc;
rom[591] = 12'hccc;
rom[592] = 12'hccc;
rom[593] = 12'hccc;
rom[594] = 12'hccc;
rom[595] = 12'hccc;
rom[596] = 12'hccc;
rom[597] = 12'hccc;
rom[598] = 12'hccc;
rom[599] = 12'h777;
rom[600] = 12'h777;
rom[601] = 12'h777;
rom[602] = 12'h777;
rom[603] = 12'h777;
rom[604] = 12'h777;
rom[605] = 12'h777;
rom[606] = 12'h777;
rom[607] = 12'h777;
rom[608] = 12'h777;
rom[609] = 12'h777;
rom[610] = 12'h777;
rom[611] = 12'h777;
rom[612] = 12'h777;
rom[613] = 12'h777;
rom[614] = 12'h777;
rom[615] = 12'h777;
rom[616] = 12'h777;
rom[617] = 12'h777;
rom[618] = 12'h777;
rom[619] = 12'h777;
rom[620] = 12'h777;
rom[621] = 12'h777;
rom[622] = 12'h777;
rom[623] = 12'h777;
rom[624] = 12'h777;
  end
endmodule

module tile_one_rom (                       //клетка с единицей
  input  wire    [13:0]     addr,
  output wire    [11:0]     word
);

  logic [11:0] rom [(25 * 25)];

  assign word = rom[addr];

  initial begin
rom[0] = 12'h777;
rom[1] = 12'h777;
rom[2] = 12'h777;
rom[3] = 12'h777;
rom[4] = 12'h777;
rom[5] = 12'h777;
rom[6] = 12'h777;
rom[7] = 12'h777;
rom[8] = 12'h777;
rom[9] = 12'h777;
rom[10] = 12'h777;
rom[11] = 12'h777;
rom[12] = 12'h777;
rom[13] = 12'h777;
rom[14] = 12'h777;
rom[15] = 12'h777;
rom[16] = 12'h777;
rom[17] = 12'h777;
rom[18] = 12'h777;
rom[19] = 12'h777;
rom[20] = 12'h777;
rom[21] = 12'h777;
rom[22] = 12'h777;
rom[23] = 12'h777;
rom[24] = 12'h777;
rom[25] = 12'h777;
rom[26] = 12'hccc;
rom[27] = 12'hccc;
rom[28] = 12'hccc;
rom[29] = 12'hccc;
rom[30] = 12'hccc;
rom[31] = 12'hccc;
rom[32] = 12'hccc;
rom[33] = 12'hccc;
rom[34] = 12'hccc;
rom[35] = 12'hccc;
rom[36] = 12'hccc;
rom[37] = 12'hccc;
rom[38] = 12'hccc;
rom[39] = 12'hccc;
rom[40] = 12'hccc;
rom[41] = 12'hccc;
rom[42] = 12'hccc;
rom[43] = 12'hccc;
rom[44] = 12'hccc;
rom[45] = 12'hccc;
rom[46] = 12'hccc;
rom[47] = 12'hccc;
rom[48] = 12'hccc;
rom[49] = 12'h777;
rom[50] = 12'h777;
rom[51] = 12'hccc;
rom[52] = 12'hccc;
rom[53] = 12'hccc;
rom[54] = 12'hccc;
rom[55] = 12'hccc;
rom[56] = 12'hccc;
rom[57] = 12'hccc;
rom[58] = 12'hccc;
rom[59] = 12'hccc;
rom[60] = 12'hccc;
rom[61] = 12'hccc;
rom[62] = 12'hccc;
rom[63] = 12'hccc;
rom[64] = 12'hccc;
rom[65] = 12'hccc;
rom[66] = 12'hccc;
rom[67] = 12'hccc;
rom[68] = 12'hccc;
rom[69] = 12'hccc;
rom[70] = 12'hccc;
rom[71] = 12'hccc;
rom[72] = 12'hccc;
rom[73] = 12'hccc;
rom[74] = 12'h777;
rom[75] = 12'h777;
rom[76] = 12'hccc;
rom[77] = 12'hccc;
rom[78] = 12'hccc;
rom[79] = 12'hccc;
rom[80] = 12'hccc;
rom[81] = 12'hccc;
rom[82] = 12'hccc;
rom[83] = 12'hccc;
rom[84] = 12'hccc;
rom[85] = 12'hccc;
rom[86] = 12'hccc;
rom[87] = 12'hccc;
rom[88] = 12'hccc;
rom[89] = 12'hccc;
rom[90] = 12'hccc;
rom[91] = 12'hccc;
rom[92] = 12'hccc;
rom[93] = 12'hccc;
rom[94] = 12'hccc;
rom[95] = 12'hccc;
rom[96] = 12'hccc;
rom[97] = 12'hccc;
rom[98] = 12'hccc;
rom[99] = 12'h777;
rom[100] = 12'h777;
rom[101] = 12'hccc;
rom[102] = 12'hccc;
rom[103] = 12'hccc;
rom[104] = 12'hccc;
rom[105] = 12'hccc;
rom[106] = 12'hccc;
rom[107] = 12'hccc;
rom[108] = 12'hccc;
rom[109] = 12'hccc;
rom[110] = 12'hccc;
rom[111] = 12'hccc;
rom[112] = 12'hccc;
rom[113] = 12'hccc;
rom[114] = 12'hccc;
rom[115] = 12'hccc;
rom[116] = 12'hccc;
rom[117] = 12'hccc;
rom[118] = 12'hccc;
rom[119] = 12'hccc;
rom[120] = 12'hccc;
rom[121] = 12'hccc;
rom[122] = 12'hccc;
rom[123] = 12'hccc;
rom[124] = 12'h777;
rom[125] = 12'h777;
rom[126] = 12'hccc;
rom[127] = 12'hccc;
rom[128] = 12'hccc;
rom[129] = 12'hccc;
rom[130] = 12'hccc;
rom[131] = 12'hccc;
rom[132] = 12'hccc;
rom[133] = 12'hccc;
rom[134] = 12'hccc;
rom[135] = 12'hccc;
rom[136] = 12'hccc;
rom[137] = 12'hccc;
rom[138] = 12'hccc;
rom[139] = 12'hccc;
rom[140] = 12'hccc;
rom[141] = 12'hccc;
rom[142] = 12'hccc;
rom[143] = 12'hccc;
rom[144] = 12'hccc;
rom[145] = 12'hccc;
rom[146] = 12'hccc;
rom[147] = 12'hccc;
rom[148] = 12'hccc;
rom[149] = 12'h777;
rom[150] = 12'h777;
rom[151] = 12'hccc;
rom[152] = 12'hccc;
rom[153] = 12'hccc;
rom[154] = 12'hccc;
rom[155] = 12'hccc;
rom[156] = 12'hccc;
rom[157] = 12'hccc;
rom[158] = 12'hccc;
rom[159] = 12'hccc;
rom[160] = 12'hccc;
rom[161] = 12'hccc;
rom[162] = 12'hccc;
rom[163] = 12'hccc;
rom[164] = 12'hccc;
rom[165] = 12'hccc;
rom[166] = 12'hccc;
rom[167] = 12'hccc;
rom[168] = 12'hccc;
rom[169] = 12'hccc;
rom[170] = 12'hccc;
rom[171] = 12'hccc;
rom[172] = 12'hccc;
rom[173] = 12'hccc;
rom[174] = 12'h777;
rom[175] = 12'h777;
rom[176] = 12'hccc;
rom[177] = 12'hccc;
rom[178] = 12'hccc;
rom[179] = 12'hccc;
rom[180] = 12'hccc;
rom[181] = 12'hccc;
rom[182] = 12'hccc;
rom[183] = 12'hccc;
rom[184] = 12'h070;
rom[185] = 12'h070;
rom[186] = 12'h070;
rom[187] = 12'h070;
rom[188] = 12'h070;
rom[189] = 12'h070;
rom[190] = 12'h070;
rom[191] = 12'h070;
rom[192] = 12'hccc;
rom[193] = 12'hccc;
rom[194] = 12'hccc;
rom[195] = 12'hccc;
rom[196] = 12'hccc;
rom[197] = 12'hccc;
rom[198] = 12'hccc;
rom[199] = 12'h777;
rom[200] = 12'h777;
rom[201] = 12'hccc;
rom[202] = 12'hccc;
rom[203] = 12'hccc;
rom[204] = 12'hccc;
rom[205] = 12'hccc;
rom[206] = 12'hccc;
rom[207] = 12'hccc;
rom[208] = 12'h070;
rom[209] = 12'h070;
rom[210] = 12'h070;
rom[211] = 12'h070;
rom[212] = 12'h070;
rom[213] = 12'h070;
rom[214] = 12'h070;
rom[215] = 12'h070;
rom[216] = 12'h070;
rom[217] = 12'h070;
rom[218] = 12'hccc;
rom[219] = 12'hccc;
rom[220] = 12'hccc;
rom[221] = 12'hccc;
rom[222] = 12'hccc;
rom[223] = 12'hccc;
rom[224] = 12'h777;
rom[225] = 12'h777;
rom[226] = 12'hccc;
rom[227] = 12'hccc;
rom[228] = 12'hccc;
rom[229] = 12'hccc;
rom[230] = 12'hccc;
rom[231] = 12'hccc;
rom[232] = 12'hccc;
rom[233] = 12'h070;
rom[234] = 12'h070;
rom[235] = 12'h070;
rom[236] = 12'hccc;
rom[237] = 12'hccc;
rom[238] = 12'hccc;
rom[239] = 12'hccc;
rom[240] = 12'h070;
rom[241] = 12'h070;
rom[242] = 12'h070;
rom[243] = 12'hccc;
rom[244] = 12'hccc;
rom[245] = 12'hccc;
rom[246] = 12'hccc;
rom[247] = 12'hccc;
rom[248] = 12'hccc;
rom[249] = 12'h777;
rom[250] = 12'h777;
rom[251] = 12'hccc;
rom[252] = 12'hccc;
rom[253] = 12'hccc;
rom[254] = 12'hccc;
rom[255] = 12'hccc;
rom[256] = 12'hccc;
rom[257] = 12'hccc;
rom[258] = 12'hccc;
rom[259] = 12'hccc;
rom[260] = 12'hccc;
rom[261] = 12'hccc;
rom[262] = 12'hccc;
rom[263] = 12'hccc;
rom[264] = 12'hccc;
rom[265] = 12'h070;
rom[266] = 12'h070;
rom[267] = 12'h070;
rom[268] = 12'hccc;
rom[269] = 12'hccc;
rom[270] = 12'hccc;
rom[271] = 12'hccc;
rom[272] = 12'hccc;
rom[273] = 12'hccc;
rom[274] = 12'h777;
rom[275] = 12'h777;
rom[276] = 12'hccc;
rom[277] = 12'hccc;
rom[278] = 12'hccc;
rom[279] = 12'hccc;
rom[280] = 12'hccc;
rom[281] = 12'hccc;
rom[282] = 12'hccc;
rom[283] = 12'hccc;
rom[284] = 12'hccc;
rom[285] = 12'hccc;
rom[286] = 12'hccc;
rom[287] = 12'hccc;
rom[288] = 12'h070;
rom[289] = 12'h070;
rom[290] = 12'h070;
rom[291] = 12'h070;
rom[292] = 12'hccc;
rom[293] = 12'hccc;
rom[294] = 12'hccc;
rom[295] = 12'hccc;
rom[296] = 12'hccc;
rom[297] = 12'hccc;
rom[298] = 12'hccc;
rom[299] = 12'h777;
rom[300] = 12'h777;
rom[301] = 12'hccc;
rom[302] = 12'hccc;
rom[303] = 12'hccc;
rom[304] = 12'hccc;
rom[305] = 12'hccc;
rom[306] = 12'hccc;
rom[307] = 12'hccc;
rom[308] = 12'hccc;
rom[309] = 12'hccc;
rom[310] = 12'hccc;
rom[311] = 12'h070;
rom[312] = 12'h070;
rom[313] = 12'h070;
rom[314] = 12'h070;
rom[315] = 12'h070;
rom[316] = 12'hccc;
rom[317] = 12'hccc;
rom[318] = 12'hccc;
rom[319] = 12'hccc;
rom[320] = 12'hccc;
rom[321] = 12'hccc;
rom[322] = 12'hccc;
rom[323] = 12'hccc;
rom[324] = 12'h777;
rom[325] = 12'h777;
rom[326] = 12'hccc;
rom[327] = 12'hccc;
rom[328] = 12'hccc;
rom[329] = 12'hccc;
rom[330] = 12'hccc;
rom[331] = 12'hccc;
rom[332] = 12'hccc;
rom[333] = 12'hccc;
rom[334] = 12'h070;
rom[335] = 12'h070;
rom[336] = 12'h070;
rom[337] = 12'h070;
rom[338] = 12'h070;
rom[339] = 12'hccc;
rom[340] = 12'hccc;
rom[341] = 12'hccc;
rom[342] = 12'hccc;
rom[343] = 12'hccc;
rom[344] = 12'hccc;
rom[345] = 12'hccc;
rom[346] = 12'hccc;
rom[347] = 12'hccc;
rom[348] = 12'hccc;
rom[349] = 12'h777;
rom[350] = 12'h777;
rom[351] = 12'hccc;
rom[352] = 12'hccc;
rom[353] = 12'hccc;
rom[354] = 12'hccc;
rom[355] = 12'hccc;
rom[356] = 12'hccc;
rom[357] = 12'hccc;
rom[358] = 12'h070;
rom[359] = 12'h070;
rom[360] = 12'h070;
rom[361] = 12'h070;
rom[362] = 12'hccc;
rom[363] = 12'hccc;
rom[364] = 12'hccc;
rom[365] = 12'hccc;
rom[366] = 12'hccc;
rom[367] = 12'hccc;
rom[368] = 12'hccc;
rom[369] = 12'hccc;
rom[370] = 12'hccc;
rom[371] = 12'hccc;
rom[372] = 12'hccc;
rom[373] = 12'hccc;
rom[374] = 12'h777;
rom[375] = 12'h777;
rom[376] = 12'hccc;
rom[377] = 12'hccc;
rom[378] = 12'hccc;
rom[379] = 12'hccc;
rom[380] = 12'hccc;
rom[381] = 12'hccc;
rom[382] = 12'hccc;
rom[383] = 12'h070;
rom[384] = 12'h070;
rom[385] = 12'h070;
rom[386] = 12'h070;
rom[387] = 12'h070;
rom[388] = 12'h070;
rom[389] = 12'h070;
rom[390] = 12'h070;
rom[391] = 12'h070;
rom[392] = 12'h070;
rom[393] = 12'hccc;
rom[394] = 12'hccc;
rom[395] = 12'hccc;
rom[396] = 12'hccc;
rom[397] = 12'hccc;
rom[398] = 12'hccc;
rom[399] = 12'h777;
rom[400] = 12'h777;
rom[401] = 12'hccc;
rom[402] = 12'hccc;
rom[403] = 12'hccc;
rom[404] = 12'hccc;
rom[405] = 12'hccc;
rom[406] = 12'hccc;
rom[407] = 12'hccc;
rom[408] = 12'h070;
rom[409] = 12'h070;
rom[410] = 12'h070;
rom[411] = 12'h070;
rom[412] = 12'h070;
rom[413] = 12'h070;
rom[414] = 12'h070;
rom[415] = 12'h070;
rom[416] = 12'h070;
rom[417] = 12'h070;
rom[418] = 12'hccc;
rom[419] = 12'hccc;
rom[420] = 12'hccc;
rom[421] = 12'hccc;
rom[422] = 12'hccc;
rom[423] = 12'hccc;
rom[424] = 12'h777;
rom[425] = 12'h777;
rom[426] = 12'hccc;
rom[427] = 12'hccc;
rom[428] = 12'hccc;
rom[429] = 12'hccc;
rom[430] = 12'hccc;
rom[431] = 12'hccc;
rom[432] = 12'hccc;
rom[433] = 12'hccc;
rom[434] = 12'hccc;
rom[435] = 12'hccc;
rom[436] = 12'hccc;
rom[437] = 12'hccc;
rom[438] = 12'hccc;
rom[439] = 12'hccc;
rom[440] = 12'hbbb;
rom[441] = 12'hccc;
rom[442] = 12'hccc;
rom[443] = 12'hccc;
rom[444] = 12'hccc;
rom[445] = 12'hccc;
rom[446] = 12'hccc;
rom[447] = 12'hccc;
rom[448] = 12'hccc;
rom[449] = 12'h777;
rom[450] = 12'h777;
rom[451] = 12'hccc;
rom[452] = 12'hccc;
rom[453] = 12'hccc;
rom[454] = 12'hccc;
rom[455] = 12'hccc;
rom[456] = 12'hccc;
rom[457] = 12'hccc;
rom[458] = 12'hccc;
rom[459] = 12'hccc;
rom[460] = 12'hccc;
rom[461] = 12'hccc;
rom[462] = 12'hccc;
rom[463] = 12'hccc;
rom[464] = 12'hccc;
rom[465] = 12'hbbb;
rom[466] = 12'hccc;
rom[467] = 12'hccc;
rom[468] = 12'hccc;
rom[469] = 12'hccc;
rom[470] = 12'hccc;
rom[471] = 12'hccc;
rom[472] = 12'hccc;
rom[473] = 12'hccc;
rom[474] = 12'h777;
rom[475] = 12'h777;
rom[476] = 12'hccc;
rom[477] = 12'hccc;
rom[478] = 12'hccc;
rom[479] = 12'hccc;
rom[480] = 12'hccc;
rom[481] = 12'hccc;
rom[482] = 12'hccc;
rom[483] = 12'hccc;
rom[484] = 12'hccc;
rom[485] = 12'hccc;
rom[486] = 12'hccc;
rom[487] = 12'hccc;
rom[488] = 12'hccc;
rom[489] = 12'hccc;
rom[490] = 12'hccc;
rom[491] = 12'hccc;
rom[492] = 12'hccc;
rom[493] = 12'hccc;
rom[494] = 12'hccc;
rom[495] = 12'hccc;
rom[496] = 12'hccc;
rom[497] = 12'hccc;
rom[498] = 12'hccc;
rom[499] = 12'h777;
rom[500] = 12'h777;
rom[501] = 12'hccc;
rom[502] = 12'hccc;
rom[503] = 12'hccc;
rom[504] = 12'hccc;
rom[505] = 12'hccc;
rom[506] = 12'hccc;
rom[507] = 12'hccc;
rom[508] = 12'hccc;
rom[509] = 12'hccc;
rom[510] = 12'hccc;
rom[511] = 12'hccc;
rom[512] = 12'hccc;
rom[513] = 12'hccc;
rom[514] = 12'hccc;
rom[515] = 12'hccc;
rom[516] = 12'hccc;
rom[517] = 12'hccc;
rom[518] = 12'hccc;
rom[519] = 12'hccc;
rom[520] = 12'hccc;
rom[521] = 12'hccc;
rom[522] = 12'hccc;
rom[523] = 12'hccc;
rom[524] = 12'h777;
rom[525] = 12'h777;
rom[526] = 12'hccc;
rom[527] = 12'hccc;
rom[528] = 12'hccc;
rom[529] = 12'hccc;
rom[530] = 12'hccc;
rom[531] = 12'hccc;
rom[532] = 12'hccc;
rom[533] = 12'hccc;
rom[534] = 12'hccc;
rom[535] = 12'hccc;
rom[536] = 12'hccc;
rom[537] = 12'hccc;
rom[538] = 12'hccc;
rom[539] = 12'hccc;
rom[540] = 12'hccc;
rom[541] = 12'hccc;
rom[542] = 12'hccc;
rom[543] = 12'hccc;
rom[544] = 12'hccc;
rom[545] = 12'hccc;
rom[546] = 12'hccc;
rom[547] = 12'hccc;
rom[548] = 12'hccc;
rom[549] = 12'h777;
rom[550] = 12'h777;
rom[551] = 12'hccc;
rom[552] = 12'hccc;
rom[553] = 12'hccc;
rom[554] = 12'hccc;
rom[555] = 12'hccc;
rom[556] = 12'hccc;
rom[557] = 12'hccc;
rom[558] = 12'hccc;
rom[559] = 12'hccc;
rom[560] = 12'hccc;
rom[561] = 12'hccc;
rom[562] = 12'hccc;
rom[563] = 12'hccc;
rom[564] = 12'hccc;
rom[565] = 12'hccc;
rom[566] = 12'hccc;
rom[567] = 12'hccc;
rom[568] = 12'hccc;
rom[569] = 12'hccc;
rom[570] = 12'hccc;
rom[571] = 12'hccc;
rom[572] = 12'hccc;
rom[573] = 12'hccc;
rom[574] = 12'h777;
rom[575] = 12'h777;
rom[576] = 12'hccc;
rom[577] = 12'hccc;
rom[578] = 12'hccc;
rom[579] = 12'hccc;
rom[580] = 12'hccc;
rom[581] = 12'hccc;
rom[582] = 12'hccc;
rom[583] = 12'hccc;
rom[584] = 12'hccc;
rom[585] = 12'hccc;
rom[586] = 12'hccc;
rom[587] = 12'hccc;
rom[588] = 12'hccc;
rom[589] = 12'hccc;
rom[590] = 12'hccc;
rom[591] = 12'hccc;
rom[592] = 12'hccc;
rom[593] = 12'hccc;
rom[594] = 12'hccc;
rom[595] = 12'hccc;
rom[596] = 12'hccc;
rom[597] = 12'hccc;
rom[598] = 12'hccc;
rom[599] = 12'h777;
rom[600] = 12'h777;
rom[601] = 12'h777;
rom[602] = 12'h777;
rom[603] = 12'h777;
rom[604] = 12'h777;
rom[605] = 12'h777;
rom[606] = 12'h777;
rom[607] = 12'h777;
rom[608] = 12'h777;
rom[609] = 12'h777;
rom[610] = 12'h777;
rom[611] = 12'h777;
rom[612] = 12'h777;
rom[613] = 12'h777;
rom[614] = 12'h777;
rom[615] = 12'h777;
rom[616] = 12'h777;
rom[617] = 12'h777;
rom[618] = 12'h777;
rom[619] = 12'h777;
rom[620] = 12'h777;
rom[621] = 12'h777;
rom[622] = 12'h777;
rom[623] = 12'h777;
rom[624] = 12'h777;
  end
endmodule

module tile_tree_rom (                       //клетка с тройкой
  input  wire    [13:0]     addr,
  output wire    [11:0]     word
);

  logic [11:0] rom [(25 * 25)];

  assign word = rom[addr];

  initial begin
rom[0] = 12'h777;
rom[1] = 12'h777;
rom[2] = 12'h777;
rom[3] = 12'h777;
rom[4] = 12'h777;
rom[5] = 12'h777;
rom[6] = 12'h777;
rom[7] = 12'h777;
rom[8] = 12'h777;
rom[9] = 12'h777;
rom[10] = 12'h777;
rom[11] = 12'h777;
rom[12] = 12'h777;
rom[13] = 12'h777;
rom[14] = 12'h777;
rom[15] = 12'h777;
rom[16] = 12'h777;
rom[17] = 12'h777;
rom[18] = 12'h777;
rom[19] = 12'h777;
rom[20] = 12'h777;
rom[21] = 12'h777;
rom[22] = 12'h777;
rom[23] = 12'h777;
rom[24] = 12'h777;
rom[25] = 12'h777;
rom[26] = 12'hccc;
rom[27] = 12'hccc;
rom[28] = 12'hccc;
rom[29] = 12'hccc;
rom[30] = 12'hccc;
rom[31] = 12'hccc;
rom[32] = 12'hccc;
rom[33] = 12'hccc;
rom[34] = 12'hccc;
rom[35] = 12'hccc;
rom[36] = 12'hccc;
rom[37] = 12'hccc;
rom[38] = 12'hccc;
rom[39] = 12'hccc;
rom[40] = 12'hccc;
rom[41] = 12'hccc;
rom[42] = 12'hccc;
rom[43] = 12'hccc;
rom[44] = 12'hccc;
rom[45] = 12'hccc;
rom[46] = 12'hccc;
rom[47] = 12'hccc;
rom[48] = 12'hccc;
rom[49] = 12'h777;
rom[50] = 12'h777;
rom[51] = 12'hccc;
rom[52] = 12'hccc;
rom[53] = 12'hccc;
rom[54] = 12'hccc;
rom[55] = 12'hccc;
rom[56] = 12'hccc;
rom[57] = 12'hccc;
rom[58] = 12'hccc;
rom[59] = 12'hccc;
rom[60] = 12'hccc;
rom[61] = 12'hccc;
rom[62] = 12'hccc;
rom[63] = 12'hccc;
rom[64] = 12'hccc;
rom[65] = 12'hccc;
rom[66] = 12'hccc;
rom[67] = 12'hccc;
rom[68] = 12'hccc;
rom[69] = 12'hccc;
rom[70] = 12'hccc;
rom[71] = 12'hccc;
rom[72] = 12'hccc;
rom[73] = 12'hccc;
rom[74] = 12'h777;
rom[75] = 12'h777;
rom[76] = 12'hccc;
rom[77] = 12'hccc;
rom[78] = 12'hccc;
rom[79] = 12'hccc;
rom[80] = 12'hccc;
rom[81] = 12'hccc;
rom[82] = 12'hccc;
rom[83] = 12'hccc;
rom[84] = 12'hccc;
rom[85] = 12'hccc;
rom[86] = 12'hccc;
rom[87] = 12'hccc;
rom[88] = 12'hccc;
rom[89] = 12'hccc;
rom[90] = 12'hccc;
rom[91] = 12'hccc;
rom[92] = 12'hccc;
rom[93] = 12'hccc;
rom[94] = 12'hccc;
rom[95] = 12'hccc;
rom[96] = 12'hccc;
rom[97] = 12'hccc;
rom[98] = 12'hccc;
rom[99] = 12'h777;
rom[100] = 12'h777;
rom[101] = 12'hccc;
rom[102] = 12'hccc;
rom[103] = 12'hccc;
rom[104] = 12'hccc;
rom[105] = 12'hccc;
rom[106] = 12'hccc;
rom[107] = 12'hccc;
rom[108] = 12'hccc;
rom[109] = 12'hccc;
rom[110] = 12'hccc;
rom[111] = 12'hccc;
rom[112] = 12'hccc;
rom[113] = 12'hccc;
rom[114] = 12'hccc;
rom[115] = 12'hccc;
rom[116] = 12'hccc;
rom[117] = 12'hccc;
rom[118] = 12'hccc;
rom[119] = 12'hccc;
rom[120] = 12'hccc;
rom[121] = 12'hccc;
rom[122] = 12'hccc;
rom[123] = 12'hccc;
rom[124] = 12'h777;
rom[125] = 12'h777;
rom[126] = 12'hccc;
rom[127] = 12'hccc;
rom[128] = 12'hccc;
rom[129] = 12'hccc;
rom[130] = 12'hccc;
rom[131] = 12'hccc;
rom[132] = 12'hccc;
rom[133] = 12'hccc;
rom[134] = 12'hccc;
rom[135] = 12'hccc;
rom[136] = 12'hccc;
rom[137] = 12'hccc;
rom[138] = 12'hccc;
rom[139] = 12'hccc;
rom[140] = 12'hccc;
rom[141] = 12'hccc;
rom[142] = 12'hccc;
rom[143] = 12'hccc;
rom[144] = 12'hccc;
rom[145] = 12'hccc;
rom[146] = 12'hccc;
rom[147] = 12'hccc;
rom[148] = 12'hccc;
rom[149] = 12'h777;
rom[150] = 12'h777;
rom[151] = 12'hccc;
rom[152] = 12'hccc;
rom[153] = 12'hccc;
rom[154] = 12'hccc;
rom[155] = 12'hccc;
rom[156] = 12'hccc;
rom[157] = 12'hccc;
rom[158] = 12'hccc;
rom[159] = 12'hccc;
rom[160] = 12'hccc;
rom[161] = 12'hccc;
rom[162] = 12'hccc;
rom[163] = 12'hccc;
rom[164] = 12'hccc;
rom[165] = 12'hccc;
rom[166] = 12'hccc;
rom[167] = 12'hccc;
rom[168] = 12'hccc;
rom[169] = 12'hccc;
rom[170] = 12'hccc;
rom[171] = 12'hccc;
rom[172] = 12'hccc;
rom[173] = 12'hccc;
rom[174] = 12'h777;
rom[175] = 12'h777;
rom[176] = 12'hccc;
rom[177] = 12'hccc;
rom[178] = 12'hccc;
rom[179] = 12'hccc;
rom[180] = 12'hccc;
rom[181] = 12'hccc;
rom[182] = 12'hccc;
rom[183] = 12'h00f;
rom[184] = 12'h00f;
rom[185] = 12'h00f;
rom[186] = 12'h00f;
rom[187] = 12'h00f;
rom[188] = 12'h00f;
rom[189] = 12'h00f;
rom[190] = 12'h00f;
rom[191] = 12'h00f;
rom[192] = 12'hccc;
rom[193] = 12'hccc;
rom[194] = 12'hccc;
rom[195] = 12'hccc;
rom[196] = 12'hccc;
rom[197] = 12'hccc;
rom[198] = 12'hccc;
rom[199] = 12'h777;
rom[200] = 12'h777;
rom[201] = 12'hccc;
rom[202] = 12'hccc;
rom[203] = 12'hccc;
rom[204] = 12'hccc;
rom[205] = 12'hccc;
rom[206] = 12'hccc;
rom[207] = 12'hccc;
rom[208] = 12'h00f;
rom[209] = 12'h00f;
rom[210] = 12'h00f;
rom[211] = 12'h00f;
rom[212] = 12'h00f;
rom[213] = 12'h00f;
rom[214] = 12'h00f;
rom[215] = 12'h00f;
rom[216] = 12'h00f;
rom[217] = 12'h00f;
rom[218] = 12'hccc;
rom[219] = 12'hccc;
rom[220] = 12'hccc;
rom[221] = 12'hccc;
rom[222] = 12'hccc;
rom[223] = 12'hccc;
rom[224] = 12'h777;
rom[225] = 12'h777;
rom[226] = 12'hccc;
rom[227] = 12'hccc;
rom[228] = 12'hccc;
rom[229] = 12'hccc;
rom[230] = 12'hccc;
rom[231] = 12'hccc;
rom[232] = 12'hccc;
rom[233] = 12'hccc;
rom[234] = 12'hccc;
rom[235] = 12'hccc;
rom[236] = 12'hccc;
rom[237] = 12'hccc;
rom[238] = 12'hccc;
rom[239] = 12'hccc;
rom[240] = 12'h00f;
rom[241] = 12'h00f;
rom[242] = 12'h00f;
rom[243] = 12'hccc;
rom[244] = 12'hccc;
rom[245] = 12'hccc;
rom[246] = 12'hccc;
rom[247] = 12'hccc;
rom[248] = 12'hccc;
rom[249] = 12'h777;
rom[250] = 12'h777;
rom[251] = 12'hccc;
rom[252] = 12'hccc;
rom[253] = 12'hccc;
rom[254] = 12'hccc;
rom[255] = 12'hccc;
rom[256] = 12'hccc;
rom[257] = 12'hccc;
rom[258] = 12'hccc;
rom[259] = 12'hccc;
rom[260] = 12'hccc;
rom[261] = 12'hccc;
rom[262] = 12'hccc;
rom[263] = 12'hccc;
rom[264] = 12'hccc;
rom[265] = 12'h00f;
rom[266] = 12'h00f;
rom[267] = 12'h00f;
rom[268] = 12'hccc;
rom[269] = 12'hccc;
rom[270] = 12'hccc;
rom[271] = 12'hccc;
rom[272] = 12'hccc;
rom[273] = 12'hccc;
rom[274] = 12'h777;
rom[275] = 12'h777;
rom[276] = 12'hccc;
rom[277] = 12'hccc;
rom[278] = 12'hccc;
rom[279] = 12'hccc;
rom[280] = 12'hccc;
rom[281] = 12'hccc;
rom[282] = 12'hccc;
rom[283] = 12'hccc;
rom[284] = 12'hccc;
rom[285] = 12'hccc;
rom[286] = 12'h00f;
rom[287] = 12'h00f;
rom[288] = 12'h00f;
rom[289] = 12'h00f;
rom[290] = 12'h00f;
rom[291] = 12'h00f;
rom[292] = 12'hccc;
rom[293] = 12'hccc;
rom[294] = 12'hccc;
rom[295] = 12'hccc;
rom[296] = 12'hccc;
rom[297] = 12'hccc;
rom[298] = 12'hccc;
rom[299] = 12'h777;
rom[300] = 12'h777;
rom[301] = 12'hccc;
rom[302] = 12'hccc;
rom[303] = 12'hccc;
rom[304] = 12'hccc;
rom[305] = 12'hccc;
rom[306] = 12'hccc;
rom[307] = 12'hccc;
rom[308] = 12'hccc;
rom[309] = 12'hccc;
rom[310] = 12'hccc;
rom[311] = 12'h00f;
rom[312] = 12'h00f;
rom[313] = 12'h00f;
rom[314] = 12'h00f;
rom[315] = 12'h00f;
rom[316] = 12'h00f;
rom[317] = 12'hccc;
rom[318] = 12'hccc;
rom[319] = 12'hccc;
rom[320] = 12'hccc;
rom[321] = 12'hccc;
rom[322] = 12'hccc;
rom[323] = 12'hccc;
rom[324] = 12'h777;
rom[325] = 12'h777;
rom[326] = 12'hccc;
rom[327] = 12'hccc;
rom[328] = 12'hccc;
rom[329] = 12'hccc;
rom[330] = 12'hccc;
rom[331] = 12'hccc;
rom[332] = 12'hccc;
rom[333] = 12'hccc;
rom[334] = 12'hccc;
rom[335] = 12'hccc;
rom[336] = 12'hccc;
rom[337] = 12'hccc;
rom[338] = 12'hccc;
rom[339] = 12'hccc;
rom[340] = 12'h00f;
rom[341] = 12'h00f;
rom[342] = 12'h00f;
rom[343] = 12'hccc;
rom[344] = 12'hccc;
rom[345] = 12'hccc;
rom[346] = 12'hccc;
rom[347] = 12'hccc;
rom[348] = 12'hccc;
rom[349] = 12'h777;
rom[350] = 12'h777;
rom[351] = 12'hccc;
rom[352] = 12'hccc;
rom[353] = 12'hccc;
rom[354] = 12'hccc;
rom[355] = 12'hccc;
rom[356] = 12'hccc;
rom[357] = 12'hccc;
rom[358] = 12'hccc;
rom[359] = 12'hccc;
rom[360] = 12'hccc;
rom[361] = 12'hccc;
rom[362] = 12'hccc;
rom[363] = 12'hccc;
rom[364] = 12'hccc;
rom[365] = 12'h00f;
rom[366] = 12'h00f;
rom[367] = 12'h00f;
rom[368] = 12'hccc;
rom[369] = 12'hccc;
rom[370] = 12'hccc;
rom[371] = 12'hccc;
rom[372] = 12'hccc;
rom[373] = 12'hccc;
rom[374] = 12'h777;
rom[375] = 12'h777;
rom[376] = 12'hccc;
rom[377] = 12'hccc;
rom[378] = 12'hccc;
rom[379] = 12'hccc;
rom[380] = 12'hccc;
rom[381] = 12'hccc;
rom[382] = 12'hccc;
rom[383] = 12'h00f;
rom[384] = 12'h00f;
rom[385] = 12'h00f;
rom[386] = 12'h00f;
rom[387] = 12'h00f;
rom[388] = 12'h00f;
rom[389] = 12'h00f;
rom[390] = 12'h00f;
rom[391] = 12'h00f;
rom[392] = 12'h00f;
rom[393] = 12'hccc;
rom[394] = 12'hccc;
rom[395] = 12'hccc;
rom[396] = 12'hccc;
rom[397] = 12'hccc;
rom[398] = 12'hccc;
rom[399] = 12'h777;
rom[400] = 12'h777;
rom[401] = 12'hccc;
rom[402] = 12'hccc;
rom[403] = 12'hccc;
rom[404] = 12'hccc;
rom[405] = 12'hccc;
rom[406] = 12'hccc;
rom[407] = 12'hccc;
rom[408] = 12'h00f;
rom[409] = 12'h00f;
rom[410] = 12'h00f;
rom[411] = 12'h00f;
rom[412] = 12'h00f;
rom[413] = 12'h00f;
rom[414] = 12'h00f;
rom[415] = 12'h00f;
rom[416] = 12'h00f;
rom[417] = 12'hccc;
rom[418] = 12'hccc;
rom[419] = 12'hccc;
rom[420] = 12'hccc;
rom[421] = 12'hccc;
rom[422] = 12'hccc;
rom[423] = 12'hccc;
rom[424] = 12'h777;
rom[425] = 12'h777;
rom[426] = 12'hccc;
rom[427] = 12'hccc;
rom[428] = 12'hccc;
rom[429] = 12'hccc;
rom[430] = 12'hccc;
rom[431] = 12'hccc;
rom[432] = 12'hccc;
rom[433] = 12'hccc;
rom[434] = 12'hccc;
rom[435] = 12'hccc;
rom[436] = 12'hccc;
rom[437] = 12'hccc;
rom[438] = 12'hccc;
rom[439] = 12'hccc;
rom[440] = 12'hbbb;
rom[441] = 12'hccc;
rom[442] = 12'hccc;
rom[443] = 12'hccc;
rom[444] = 12'hccc;
rom[445] = 12'hccc;
rom[446] = 12'hccc;
rom[447] = 12'hccc;
rom[448] = 12'hccc;
rom[449] = 12'h777;
rom[450] = 12'h777;
rom[451] = 12'hccc;
rom[452] = 12'hccc;
rom[453] = 12'hccc;
rom[454] = 12'hccc;
rom[455] = 12'hccc;
rom[456] = 12'hccc;
rom[457] = 12'hccc;
rom[458] = 12'hccc;
rom[459] = 12'hccc;
rom[460] = 12'hccc;
rom[461] = 12'hccc;
rom[462] = 12'hccc;
rom[463] = 12'hccc;
rom[464] = 12'hccc;
rom[465] = 12'hbbb;
rom[466] = 12'hccc;
rom[467] = 12'hccc;
rom[468] = 12'hccc;
rom[469] = 12'hccc;
rom[470] = 12'hccc;
rom[471] = 12'hccc;
rom[472] = 12'hccc;
rom[473] = 12'hccc;
rom[474] = 12'h777;
rom[475] = 12'h777;
rom[476] = 12'hccc;
rom[477] = 12'hccc;
rom[478] = 12'hccc;
rom[479] = 12'hccc;
rom[480] = 12'hccc;
rom[481] = 12'hccc;
rom[482] = 12'hccc;
rom[483] = 12'hccc;
rom[484] = 12'hccc;
rom[485] = 12'hccc;
rom[486] = 12'hccc;
rom[487] = 12'hccc;
rom[488] = 12'hccc;
rom[489] = 12'hccc;
rom[490] = 12'hccc;
rom[491] = 12'hccc;
rom[492] = 12'hccc;
rom[493] = 12'hccc;
rom[494] = 12'hccc;
rom[495] = 12'hccc;
rom[496] = 12'hccc;
rom[497] = 12'hccc;
rom[498] = 12'hccc;
rom[499] = 12'h777;
rom[500] = 12'h777;
rom[501] = 12'hccc;
rom[502] = 12'hccc;
rom[503] = 12'hccc;
rom[504] = 12'hccc;
rom[505] = 12'hccc;
rom[506] = 12'hccc;
rom[507] = 12'hccc;
rom[508] = 12'hccc;
rom[509] = 12'hccc;
rom[510] = 12'hccc;
rom[511] = 12'hccc;
rom[512] = 12'hccc;
rom[513] = 12'hccc;
rom[514] = 12'hccc;
rom[515] = 12'hccc;
rom[516] = 12'hccc;
rom[517] = 12'hccc;
rom[518] = 12'hccc;
rom[519] = 12'hccc;
rom[520] = 12'hccc;
rom[521] = 12'hccc;
rom[522] = 12'hccc;
rom[523] = 12'hccc;
rom[524] = 12'h777;
rom[525] = 12'h777;
rom[526] = 12'hccc;
rom[527] = 12'hccc;
rom[528] = 12'hccc;
rom[529] = 12'hccc;
rom[530] = 12'hccc;
rom[531] = 12'hccc;
rom[532] = 12'hccc;
rom[533] = 12'hccc;
rom[534] = 12'hccc;
rom[535] = 12'hccc;
rom[536] = 12'hccc;
rom[537] = 12'hccc;
rom[538] = 12'hccc;
rom[539] = 12'hccc;
rom[540] = 12'hccc;
rom[541] = 12'hccc;
rom[542] = 12'hccc;
rom[543] = 12'hccc;
rom[544] = 12'hccc;
rom[545] = 12'hccc;
rom[546] = 12'hccc;
rom[547] = 12'hccc;
rom[548] = 12'hccc;
rom[549] = 12'h777;
rom[550] = 12'h777;
rom[551] = 12'hccc;
rom[552] = 12'hccc;
rom[553] = 12'hccc;
rom[554] = 12'hccc;
rom[555] = 12'hccc;
rom[556] = 12'hccc;
rom[557] = 12'hccc;
rom[558] = 12'hccc;
rom[559] = 12'hccc;
rom[560] = 12'hccc;
rom[561] = 12'hccc;
rom[562] = 12'hccc;
rom[563] = 12'hccc;
rom[564] = 12'hccc;
rom[565] = 12'hccc;
rom[566] = 12'hccc;
rom[567] = 12'hccc;
rom[568] = 12'hccc;
rom[569] = 12'hccc;
rom[570] = 12'hccc;
rom[571] = 12'hccc;
rom[572] = 12'hccc;
rom[573] = 12'hccc;
rom[574] = 12'h777;
rom[575] = 12'h777;
rom[576] = 12'hccc;
rom[577] = 12'hccc;
rom[578] = 12'hccc;
rom[579] = 12'hccc;
rom[580] = 12'hccc;
rom[581] = 12'hccc;
rom[582] = 12'hccc;
rom[583] = 12'hccc;
rom[584] = 12'hccc;
rom[585] = 12'hccc;
rom[586] = 12'hccc;
rom[587] = 12'hccc;
rom[588] = 12'hccc;
rom[589] = 12'hccc;
rom[590] = 12'hccc;
rom[591] = 12'hccc;
rom[592] = 12'hccc;
rom[593] = 12'hccc;
rom[594] = 12'hccc;
rom[595] = 12'hccc;
rom[596] = 12'hccc;
rom[597] = 12'hccc;
rom[598] = 12'hccc;
rom[599] = 12'h777;
rom[600] = 12'h777;
rom[601] = 12'h777;
rom[602] = 12'h777;
rom[603] = 12'h777;
rom[604] = 12'h777;
rom[605] = 12'h777;
rom[606] = 12'h777;
rom[607] = 12'h777;
rom[608] = 12'h777;
rom[609] = 12'h777;
rom[610] = 12'h777;
rom[611] = 12'h777;
rom[612] = 12'h777;
rom[613] = 12'h777;
rom[614] = 12'h777;
rom[615] = 12'h777;
rom[616] = 12'h777;
rom[617] = 12'h777;
rom[618] = 12'h777;
rom[619] = 12'h777;
rom[620] = 12'h777;
rom[621] = 12'h777;
rom[622] = 12'h777;
rom[623] = 12'h777;
rom[624] = 12'h777;
  end
endmodule

module tile_four_rom (                       //клетка с четвёркой
  input  wire    [13:0]     addr,
  output wire    [11:0]     word
);

  logic [11:0] rom [(25 * 25)];

  assign word = rom[addr];

  initial begin
rom[0] = 12'h777;
rom[1] = 12'h777;
rom[2] = 12'h777;
rom[3] = 12'h777;
rom[4] = 12'h777;
rom[5] = 12'h777;
rom[6] = 12'h777;
rom[7] = 12'h777;
rom[8] = 12'h777;
rom[9] = 12'h777;
rom[10] = 12'h777;
rom[11] = 12'h777;
rom[12] = 12'h777;
rom[13] = 12'h777;
rom[14] = 12'h777;
rom[15] = 12'h777;
rom[16] = 12'h777;
rom[17] = 12'h777;
rom[18] = 12'h777;
rom[19] = 12'h777;
rom[20] = 12'h777;
rom[21] = 12'h777;
rom[22] = 12'h777;
rom[23] = 12'h777;
rom[24] = 12'h777;
rom[25] = 12'h777;
rom[26] = 12'hccc;
rom[27] = 12'hccc;
rom[28] = 12'hccc;
rom[29] = 12'hccc;
rom[30] = 12'hccc;
rom[31] = 12'hccc;
rom[32] = 12'hccc;
rom[33] = 12'hccc;
rom[34] = 12'hccc;
rom[35] = 12'hccc;
rom[36] = 12'hccc;
rom[37] = 12'hccc;
rom[38] = 12'hccc;
rom[39] = 12'hccc;
rom[40] = 12'hccc;
rom[41] = 12'hccc;
rom[42] = 12'hccc;
rom[43] = 12'hccc;
rom[44] = 12'hccc;
rom[45] = 12'hccc;
rom[46] = 12'hccc;
rom[47] = 12'hccc;
rom[48] = 12'hccc;
rom[49] = 12'h777;
rom[50] = 12'h777;
rom[51] = 12'hccc;
rom[52] = 12'hccc;
rom[53] = 12'hccc;
rom[54] = 12'hccc;
rom[55] = 12'hccc;
rom[56] = 12'hccc;
rom[57] = 12'hccc;
rom[58] = 12'hccc;
rom[59] = 12'hccc;
rom[60] = 12'hccc;
rom[61] = 12'hccc;
rom[62] = 12'hccc;
rom[63] = 12'hccc;
rom[64] = 12'hccc;
rom[65] = 12'hccc;
rom[66] = 12'hccc;
rom[67] = 12'hccc;
rom[68] = 12'hccc;
rom[69] = 12'hccc;
rom[70] = 12'hccc;
rom[71] = 12'hccc;
rom[72] = 12'hccc;
rom[73] = 12'hccc;
rom[74] = 12'h777;
rom[75] = 12'h777;
rom[76] = 12'hccc;
rom[77] = 12'hccc;
rom[78] = 12'hccc;
rom[79] = 12'hccc;
rom[80] = 12'hccc;
rom[81] = 12'hccc;
rom[82] = 12'hccc;
rom[83] = 12'hccc;
rom[84] = 12'hccc;
rom[85] = 12'hccc;
rom[86] = 12'hccc;
rom[87] = 12'hccc;
rom[88] = 12'hccc;
rom[89] = 12'hccc;
rom[90] = 12'hccc;
rom[91] = 12'hccc;
rom[92] = 12'hccc;
rom[93] = 12'hccc;
rom[94] = 12'hccc;
rom[95] = 12'hccc;
rom[96] = 12'hccc;
rom[97] = 12'hccc;
rom[98] = 12'hccc;
rom[99] = 12'h777;
rom[100] = 12'h777;
rom[101] = 12'hccc;
rom[102] = 12'hccc;
rom[103] = 12'hccc;
rom[104] = 12'hccc;
rom[105] = 12'hccc;
rom[106] = 12'hccc;
rom[107] = 12'hccc;
rom[108] = 12'hccc;
rom[109] = 12'hccc;
rom[110] = 12'hccc;
rom[111] = 12'hccc;
rom[112] = 12'hccc;
rom[113] = 12'hccc;
rom[114] = 12'hccc;
rom[115] = 12'hccc;
rom[116] = 12'hccc;
rom[117] = 12'hccc;
rom[118] = 12'hccc;
rom[119] = 12'hccc;
rom[120] = 12'hccc;
rom[121] = 12'hccc;
rom[122] = 12'hccc;
rom[123] = 12'hccc;
rom[124] = 12'h777;
rom[125] = 12'h777;
rom[126] = 12'hccc;
rom[127] = 12'hccc;
rom[128] = 12'hccc;
rom[129] = 12'hccc;
rom[130] = 12'hccc;
rom[131] = 12'hccc;
rom[132] = 12'hccc;
rom[133] = 12'hccc;
rom[134] = 12'hccc;
rom[135] = 12'hccc;
rom[136] = 12'hccc;
rom[137] = 12'hccc;
rom[138] = 12'hccc;
rom[139] = 12'hccc;
rom[140] = 12'hccc;
rom[141] = 12'hccc;
rom[142] = 12'hccc;
rom[143] = 12'hccc;
rom[144] = 12'hccc;
rom[145] = 12'hccc;
rom[146] = 12'hccc;
rom[147] = 12'hccc;
rom[148] = 12'hccc;
rom[149] = 12'h777;
rom[150] = 12'h777;
rom[151] = 12'hccc;
rom[152] = 12'hccc;
rom[153] = 12'hccc;
rom[154] = 12'hccc;
rom[155] = 12'hccc;
rom[156] = 12'hccc;
rom[157] = 12'hccc;
rom[158] = 12'hccc;
rom[159] = 12'hccc;
rom[160] = 12'hccc;
rom[161] = 12'hccc;
rom[162] = 12'hccc;
rom[163] = 12'hccc;
rom[164] = 12'hccc;
rom[165] = 12'hccc;
rom[166] = 12'hccc;
rom[167] = 12'hccc;
rom[168] = 12'hccc;
rom[169] = 12'hccc;
rom[170] = 12'hccc;
rom[171] = 12'hccc;
rom[172] = 12'hccc;
rom[173] = 12'hccc;
rom[174] = 12'h777;
rom[175] = 12'h777;
rom[176] = 12'hccc;
rom[177] = 12'hccc;
rom[178] = 12'hccc;
rom[179] = 12'hccc;
rom[180] = 12'hccc;
rom[181] = 12'hccc;
rom[182] = 12'hccc;
rom[183] = 12'hccc;
rom[184] = 12'h700;
rom[185] = 12'h700;
rom[186] = 12'h700;
rom[187] = 12'hccc;
rom[188] = 12'h700;
rom[189] = 12'h700;
rom[190] = 12'h700;
rom[191] = 12'hccc;
rom[192] = 12'hccc;
rom[193] = 12'hccc;
rom[194] = 12'hccc;
rom[195] = 12'hccc;
rom[196] = 12'hccc;
rom[197] = 12'hccc;
rom[198] = 12'hccc;
rom[199] = 12'h777;
rom[200] = 12'h777;
rom[201] = 12'hccc;
rom[202] = 12'hccc;
rom[203] = 12'hccc;
rom[204] = 12'hccc;
rom[205] = 12'hccc;
rom[206] = 12'hccc;
rom[207] = 12'hccc;
rom[208] = 12'hccc;
rom[209] = 12'h700;
rom[210] = 12'h700;
rom[211] = 12'h700;
rom[212] = 12'hccc;
rom[213] = 12'h700;
rom[214] = 12'h700;
rom[215] = 12'h700;
rom[216] = 12'hccc;
rom[217] = 12'hccc;
rom[218] = 12'hccc;
rom[219] = 12'hccc;
rom[220] = 12'hccc;
rom[221] = 12'hccc;
rom[222] = 12'hccc;
rom[223] = 12'hccc;
rom[224] = 12'h777;
rom[225] = 12'h777;
rom[226] = 12'hccc;
rom[227] = 12'hccc;
rom[228] = 12'hccc;
rom[229] = 12'hccc;
rom[230] = 12'hccc;
rom[231] = 12'hccc;
rom[232] = 12'hccc;
rom[233] = 12'h700;
rom[234] = 12'h700;
rom[235] = 12'h700;
rom[236] = 12'hccc;
rom[237] = 12'hccc;
rom[238] = 12'h700;
rom[239] = 12'h700;
rom[240] = 12'h700;
rom[241] = 12'hccc;
rom[242] = 12'hccc;
rom[243] = 12'hccc;
rom[244] = 12'hccc;
rom[245] = 12'hccc;
rom[246] = 12'hccc;
rom[247] = 12'hccc;
rom[248] = 12'hccc;
rom[249] = 12'h777;
rom[250] = 12'h777;
rom[251] = 12'hccc;
rom[252] = 12'hccc;
rom[253] = 12'hccc;
rom[254] = 12'hccc;
rom[255] = 12'hccc;
rom[256] = 12'hccc;
rom[257] = 12'hccc;
rom[258] = 12'h700;
rom[259] = 12'h700;
rom[260] = 12'h700;
rom[261] = 12'hccc;
rom[262] = 12'hccc;
rom[263] = 12'h700;
rom[264] = 12'h700;
rom[265] = 12'h700;
rom[266] = 12'hccc;
rom[267] = 12'hccc;
rom[268] = 12'hccc;
rom[269] = 12'hccc;
rom[270] = 12'hccc;
rom[271] = 12'hccc;
rom[272] = 12'hccc;
rom[273] = 12'hccc;
rom[274] = 12'h777;
rom[275] = 12'h777;
rom[276] = 12'hccc;
rom[277] = 12'hccc;
rom[278] = 12'hccc;
rom[279] = 12'hccc;
rom[280] = 12'hccc;
rom[281] = 12'hccc;
rom[282] = 12'h700;
rom[283] = 12'h700;
rom[284] = 12'h700;
rom[285] = 12'h700;
rom[286] = 12'h700;
rom[287] = 12'h700;
rom[288] = 12'h700;
rom[289] = 12'h700;
rom[290] = 12'h700;
rom[291] = 12'h700;
rom[292] = 12'hccc;
rom[293] = 12'hccc;
rom[294] = 12'hccc;
rom[295] = 12'hccc;
rom[296] = 12'hccc;
rom[297] = 12'hccc;
rom[298] = 12'hccc;
rom[299] = 12'h777;
rom[300] = 12'h777;
rom[301] = 12'hccc;
rom[302] = 12'hccc;
rom[303] = 12'hccc;
rom[304] = 12'hccc;
rom[305] = 12'hccc;
rom[306] = 12'hccc;
rom[307] = 12'h700;
rom[308] = 12'h700;
rom[309] = 12'h700;
rom[310] = 12'h700;
rom[311] = 12'h700;
rom[312] = 12'h700;
rom[313] = 12'h700;
rom[314] = 12'h700;
rom[315] = 12'h700;
rom[316] = 12'h700;
rom[317] = 12'hccc;
rom[318] = 12'hccc;
rom[319] = 12'hccc;
rom[320] = 12'hccc;
rom[321] = 12'hccc;
rom[322] = 12'hccc;
rom[323] = 12'hccc;
rom[324] = 12'h777;
rom[325] = 12'h777;
rom[326] = 12'hccc;
rom[327] = 12'hccc;
rom[328] = 12'hccc;
rom[329] = 12'hccc;
rom[330] = 12'hccc;
rom[331] = 12'hccc;
rom[332] = 12'hccc;
rom[333] = 12'hccc;
rom[334] = 12'hccc;
rom[335] = 12'hccc;
rom[336] = 12'hccc;
rom[337] = 12'hccc;
rom[338] = 12'h700;
rom[339] = 12'h700;
rom[340] = 12'h700;
rom[341] = 12'hccc;
rom[342] = 12'hccc;
rom[343] = 12'hccc;
rom[344] = 12'hccc;
rom[345] = 12'hccc;
rom[346] = 12'hccc;
rom[347] = 12'hccc;
rom[348] = 12'hccc;
rom[349] = 12'h777;
rom[350] = 12'h777;
rom[351] = 12'hccc;
rom[352] = 12'hccc;
rom[353] = 12'hccc;
rom[354] = 12'hccc;
rom[355] = 12'hccc;
rom[356] = 12'hccc;
rom[357] = 12'hccc;
rom[358] = 12'hccc;
rom[359] = 12'hccc;
rom[360] = 12'hccc;
rom[361] = 12'hccc;
rom[362] = 12'hccc;
rom[363] = 12'h700;
rom[364] = 12'h700;
rom[365] = 12'h700;
rom[366] = 12'hccc;
rom[367] = 12'hccc;
rom[368] = 12'hccc;
rom[369] = 12'hccc;
rom[370] = 12'hccc;
rom[371] = 12'hccc;
rom[372] = 12'hccc;
rom[373] = 12'hccc;
rom[374] = 12'h777;
rom[375] = 12'h777;
rom[376] = 12'hccc;
rom[377] = 12'hccc;
rom[378] = 12'hccc;
rom[379] = 12'hccc;
rom[380] = 12'hccc;
rom[381] = 12'hccc;
rom[382] = 12'hccc;
rom[383] = 12'hccc;
rom[384] = 12'hccc;
rom[385] = 12'hccc;
rom[386] = 12'hccc;
rom[387] = 12'hccc;
rom[388] = 12'h700;
rom[389] = 12'h700;
rom[390] = 12'h700;
rom[391] = 12'hccc;
rom[392] = 12'hccc;
rom[393] = 12'hccc;
rom[394] = 12'hccc;
rom[395] = 12'hccc;
rom[396] = 12'hccc;
rom[397] = 12'hccc;
rom[398] = 12'hccc;
rom[399] = 12'h777;
rom[400] = 12'h777;
rom[401] = 12'hccc;
rom[402] = 12'hccc;
rom[403] = 12'hccc;
rom[404] = 12'hccc;
rom[405] = 12'hccc;
rom[406] = 12'hccc;
rom[407] = 12'hccc;
rom[408] = 12'hccc;
rom[409] = 12'hccc;
rom[410] = 12'hccc;
rom[411] = 12'hccc;
rom[412] = 12'hccc;
rom[413] = 12'h700;
rom[414] = 12'h700;
rom[415] = 12'h700;
rom[416] = 12'hccc;
rom[417] = 12'hccc;
rom[418] = 12'hccc;
rom[419] = 12'hccc;
rom[420] = 12'hccc;
rom[421] = 12'hccc;
rom[422] = 12'hccc;
rom[423] = 12'hccc;
rom[424] = 12'h777;
rom[425] = 12'h777;
rom[426] = 12'hccc;
rom[427] = 12'hccc;
rom[428] = 12'hccc;
rom[429] = 12'hccc;
rom[430] = 12'hccc;
rom[431] = 12'hccc;
rom[432] = 12'hccc;
rom[433] = 12'hccc;
rom[434] = 12'hccc;
rom[435] = 12'hccc;
rom[436] = 12'hccc;
rom[437] = 12'hccc;
rom[438] = 12'hccc;
rom[439] = 12'hccc;
rom[440] = 12'hbbb;
rom[441] = 12'hccc;
rom[442] = 12'hccc;
rom[443] = 12'hccc;
rom[444] = 12'hccc;
rom[445] = 12'hccc;
rom[446] = 12'hccc;
rom[447] = 12'hccc;
rom[448] = 12'hccc;
rom[449] = 12'h777;
rom[450] = 12'h777;
rom[451] = 12'hccc;
rom[452] = 12'hccc;
rom[453] = 12'hccc;
rom[454] = 12'hccc;
rom[455] = 12'hccc;
rom[456] = 12'hccc;
rom[457] = 12'hccc;
rom[458] = 12'hccc;
rom[459] = 12'hccc;
rom[460] = 12'hccc;
rom[461] = 12'hccc;
rom[462] = 12'hccc;
rom[463] = 12'hccc;
rom[464] = 12'hccc;
rom[465] = 12'hbbb;
rom[466] = 12'hccc;
rom[467] = 12'hccc;
rom[468] = 12'hccc;
rom[469] = 12'hccc;
rom[470] = 12'hccc;
rom[471] = 12'hccc;
rom[472] = 12'hccc;
rom[473] = 12'hccc;
rom[474] = 12'h777;
rom[475] = 12'h777;
rom[476] = 12'hccc;
rom[477] = 12'hccc;
rom[478] = 12'hccc;
rom[479] = 12'hccc;
rom[480] = 12'hccc;
rom[481] = 12'hccc;
rom[482] = 12'hccc;
rom[483] = 12'hccc;
rom[484] = 12'hccc;
rom[485] = 12'hccc;
rom[486] = 12'hccc;
rom[487] = 12'hccc;
rom[488] = 12'hccc;
rom[489] = 12'hccc;
rom[490] = 12'hccc;
rom[491] = 12'hccc;
rom[492] = 12'hccc;
rom[493] = 12'hccc;
rom[494] = 12'hccc;
rom[495] = 12'hccc;
rom[496] = 12'hccc;
rom[497] = 12'hccc;
rom[498] = 12'hccc;
rom[499] = 12'h777;
rom[500] = 12'h777;
rom[501] = 12'hccc;
rom[502] = 12'hccc;
rom[503] = 12'hccc;
rom[504] = 12'hccc;
rom[505] = 12'hccc;
rom[506] = 12'hccc;
rom[507] = 12'hccc;
rom[508] = 12'hccc;
rom[509] = 12'hccc;
rom[510] = 12'hccc;
rom[511] = 12'hccc;
rom[512] = 12'hccc;
rom[513] = 12'hccc;
rom[514] = 12'hccc;
rom[515] = 12'hccc;
rom[516] = 12'hccc;
rom[517] = 12'hccc;
rom[518] = 12'hccc;
rom[519] = 12'hccc;
rom[520] = 12'hccc;
rom[521] = 12'hccc;
rom[522] = 12'hccc;
rom[523] = 12'hccc;
rom[524] = 12'h777;
rom[525] = 12'h777;
rom[526] = 12'hccc;
rom[527] = 12'hccc;
rom[528] = 12'hccc;
rom[529] = 12'hccc;
rom[530] = 12'hccc;
rom[531] = 12'hccc;
rom[532] = 12'hccc;
rom[533] = 12'hccc;
rom[534] = 12'hccc;
rom[535] = 12'hccc;
rom[536] = 12'hccc;
rom[537] = 12'hccc;
rom[538] = 12'hccc;
rom[539] = 12'hccc;
rom[540] = 12'hccc;
rom[541] = 12'hccc;
rom[542] = 12'hccc;
rom[543] = 12'hccc;
rom[544] = 12'hccc;
rom[545] = 12'hccc;
rom[546] = 12'hccc;
rom[547] = 12'hccc;
rom[548] = 12'hccc;
rom[549] = 12'h777;
rom[550] = 12'h777;
rom[551] = 12'hccc;
rom[552] = 12'hccc;
rom[553] = 12'hccc;
rom[554] = 12'hccc;
rom[555] = 12'hccc;
rom[556] = 12'hccc;
rom[557] = 12'hccc;
rom[558] = 12'hccc;
rom[559] = 12'hccc;
rom[560] = 12'hccc;
rom[561] = 12'hccc;
rom[562] = 12'hccc;
rom[563] = 12'hccc;
rom[564] = 12'hccc;
rom[565] = 12'hccc;
rom[566] = 12'hccc;
rom[567] = 12'hccc;
rom[568] = 12'hccc;
rom[569] = 12'hccc;
rom[570] = 12'hccc;
rom[571] = 12'hccc;
rom[572] = 12'hccc;
rom[573] = 12'hccc;
rom[574] = 12'h777;
rom[575] = 12'h777;
rom[576] = 12'hccc;
rom[577] = 12'hccc;
rom[578] = 12'hccc;
rom[579] = 12'hccc;
rom[580] = 12'hccc;
rom[581] = 12'hccc;
rom[582] = 12'hccc;
rom[583] = 12'hccc;
rom[584] = 12'hccc;
rom[585] = 12'hccc;
rom[586] = 12'hccc;
rom[587] = 12'hccc;
rom[588] = 12'hccc;
rom[589] = 12'hccc;
rom[590] = 12'hccc;
rom[591] = 12'hccc;
rom[592] = 12'hccc;
rom[593] = 12'hccc;
rom[594] = 12'hccc;
rom[595] = 12'hccc;
rom[596] = 12'hccc;
rom[597] = 12'hccc;
rom[598] = 12'hccc;
rom[599] = 12'h777;
rom[600] = 12'h777;
rom[601] = 12'h777;
rom[602] = 12'h777;
rom[603] = 12'h777;
rom[604] = 12'h777;
rom[605] = 12'h777;
rom[606] = 12'h777;
rom[607] = 12'h777;
rom[608] = 12'h777;
rom[609] = 12'h777;
rom[610] = 12'h777;
rom[611] = 12'h777;
rom[612] = 12'h777;
rom[613] = 12'h777;
rom[614] = 12'h777;
rom[615] = 12'h777;
rom[616] = 12'h777;
rom[617] = 12'h777;
rom[618] = 12'h777;
rom[619] = 12'h777;
rom[620] = 12'h777;
rom[621] = 12'h777;
rom[622] = 12'h777;
rom[623] = 12'h777;
rom[624] = 12'h777;
  end
endmodule

module tile_five_rom (                       //клетка с пятёркой
  input  wire    [13:0]     addr,
  output wire    [11:0]     word
);

  logic [11:0] rom [(25 * 25)];

  assign word = rom[addr];

  initial begin
rom[0] = 12'h777;
rom[1] = 12'h777;
rom[2] = 12'h777;
rom[3] = 12'h777;
rom[4] = 12'h777;
rom[5] = 12'h777;
rom[6] = 12'h777;
rom[7] = 12'h777;
rom[8] = 12'h777;
rom[9] = 12'h777;
rom[10] = 12'h777;
rom[11] = 12'h777;
rom[12] = 12'h777;
rom[13] = 12'h777;
rom[14] = 12'h777;
rom[15] = 12'h777;
rom[16] = 12'h777;
rom[17] = 12'h777;
rom[18] = 12'h777;
rom[19] = 12'h777;
rom[20] = 12'h777;
rom[21] = 12'h777;
rom[22] = 12'h777;
rom[23] = 12'h777;
rom[24] = 12'h777;
rom[25] = 12'h777;
rom[26] = 12'hccc;
rom[27] = 12'hccc;
rom[28] = 12'hccc;
rom[29] = 12'hccc;
rom[30] = 12'hccc;
rom[31] = 12'hccc;
rom[32] = 12'hccc;
rom[33] = 12'hccc;
rom[34] = 12'hccc;
rom[35] = 12'hccc;
rom[36] = 12'hccc;
rom[37] = 12'hccc;
rom[38] = 12'hccc;
rom[39] = 12'hccc;
rom[40] = 12'hccc;
rom[41] = 12'hccc;
rom[42] = 12'hccc;
rom[43] = 12'hccc;
rom[44] = 12'hccc;
rom[45] = 12'hccc;
rom[46] = 12'hccc;
rom[47] = 12'hccc;
rom[48] = 12'hccc;
rom[49] = 12'h777;
rom[50] = 12'h777;
rom[51] = 12'hccc;
rom[52] = 12'hccc;
rom[53] = 12'hccc;
rom[54] = 12'hccc;
rom[55] = 12'hccc;
rom[56] = 12'hccc;
rom[57] = 12'hccc;
rom[58] = 12'hccc;
rom[59] = 12'hccc;
rom[60] = 12'hccc;
rom[61] = 12'hccc;
rom[62] = 12'hccc;
rom[63] = 12'hccc;
rom[64] = 12'hccc;
rom[65] = 12'hccc;
rom[66] = 12'hccc;
rom[67] = 12'hccc;
rom[68] = 12'hccc;
rom[69] = 12'hccc;
rom[70] = 12'hccc;
rom[71] = 12'hccc;
rom[72] = 12'hccc;
rom[73] = 12'hccc;
rom[74] = 12'h777;
rom[75] = 12'h777;
rom[76] = 12'hccc;
rom[77] = 12'hccc;
rom[78] = 12'hccc;
rom[79] = 12'hccc;
rom[80] = 12'hccc;
rom[81] = 12'hccc;
rom[82] = 12'hccc;
rom[83] = 12'hccc;
rom[84] = 12'hccc;
rom[85] = 12'hccc;
rom[86] = 12'hccc;
rom[87] = 12'hccc;
rom[88] = 12'hccc;
rom[89] = 12'hccc;
rom[90] = 12'hccc;
rom[91] = 12'hccc;
rom[92] = 12'hccc;
rom[93] = 12'hccc;
rom[94] = 12'hccc;
rom[95] = 12'hccc;
rom[96] = 12'hccc;
rom[97] = 12'hccc;
rom[98] = 12'hccc;
rom[99] = 12'h777;
rom[100] = 12'h777;
rom[101] = 12'hccc;
rom[102] = 12'hccc;
rom[103] = 12'hccc;
rom[104] = 12'hccc;
rom[105] = 12'hccc;
rom[106] = 12'hccc;
rom[107] = 12'hccc;
rom[108] = 12'hccc;
rom[109] = 12'hccc;
rom[110] = 12'hccc;
rom[111] = 12'hccc;
rom[112] = 12'hccc;
rom[113] = 12'hccc;
rom[114] = 12'hccc;
rom[115] = 12'hccc;
rom[116] = 12'hccc;
rom[117] = 12'hccc;
rom[118] = 12'hccc;
rom[119] = 12'hccc;
rom[120] = 12'hccc;
rom[121] = 12'hccc;
rom[122] = 12'hccc;
rom[123] = 12'hccc;
rom[124] = 12'h777;
rom[125] = 12'h777;
rom[126] = 12'hccc;
rom[127] = 12'hccc;
rom[128] = 12'hccc;
rom[129] = 12'hccc;
rom[130] = 12'hccc;
rom[131] = 12'hccc;
rom[132] = 12'hccc;
rom[133] = 12'hccc;
rom[134] = 12'hccc;
rom[135] = 12'hccc;
rom[136] = 12'hccc;
rom[137] = 12'hccc;
rom[138] = 12'hccc;
rom[139] = 12'hccc;
rom[140] = 12'hccc;
rom[141] = 12'hccc;
rom[142] = 12'hccc;
rom[143] = 12'hccc;
rom[144] = 12'hccc;
rom[145] = 12'hccc;
rom[146] = 12'hccc;
rom[147] = 12'hccc;
rom[148] = 12'hccc;
rom[149] = 12'h777;
rom[150] = 12'h777;
rom[151] = 12'hccc;
rom[152] = 12'hccc;
rom[153] = 12'hccc;
rom[154] = 12'hccc;
rom[155] = 12'hccc;
rom[156] = 12'hccc;
rom[157] = 12'hccc;
rom[158] = 12'hccc;
rom[159] = 12'hccc;
rom[160] = 12'hccc;
rom[161] = 12'hccc;
rom[162] = 12'hccc;
rom[163] = 12'hccc;
rom[164] = 12'hccc;
rom[165] = 12'hccc;
rom[166] = 12'hccc;
rom[167] = 12'hccc;
rom[168] = 12'hccc;
rom[169] = 12'hccc;
rom[170] = 12'hccc;
rom[171] = 12'hccc;
rom[172] = 12'hccc;
rom[173] = 12'hccc;
rom[174] = 12'h777;
rom[175] = 12'h777;
rom[176] = 12'hccc;
rom[177] = 12'hccc;
rom[178] = 12'hccc;
rom[179] = 12'hccc;
rom[180] = 12'hccc;
rom[181] = 12'hccc;
rom[182] = 12'hccc;
rom[183] = 12'h007;
rom[184] = 12'h007;
rom[185] = 12'h007;
rom[186] = 12'h007;
rom[187] = 12'h007;
rom[188] = 12'h007;
rom[189] = 12'h007;
rom[190] = 12'h007;
rom[191] = 12'h007;
rom[192] = 12'h007;
rom[193] = 12'hccc;
rom[194] = 12'hccc;
rom[195] = 12'hccc;
rom[196] = 12'hccc;
rom[197] = 12'hccc;
rom[198] = 12'hccc;
rom[199] = 12'h777;
rom[200] = 12'h777;
rom[201] = 12'hccc;
rom[202] = 12'hccc;
rom[203] = 12'hccc;
rom[204] = 12'hccc;
rom[205] = 12'hccc;
rom[206] = 12'hccc;
rom[207] = 12'hccc;
rom[208] = 12'h007;
rom[209] = 12'h007;
rom[210] = 12'h007;
rom[211] = 12'h007;
rom[212] = 12'h007;
rom[213] = 12'h007;
rom[214] = 12'h007;
rom[215] = 12'h007;
rom[216] = 12'h007;
rom[217] = 12'h007;
rom[218] = 12'hccc;
rom[219] = 12'hccc;
rom[220] = 12'hccc;
rom[221] = 12'hccc;
rom[222] = 12'hccc;
rom[223] = 12'hccc;
rom[224] = 12'h777;
rom[225] = 12'h777;
rom[226] = 12'hccc;
rom[227] = 12'hccc;
rom[228] = 12'hccc;
rom[229] = 12'hccc;
rom[230] = 12'hccc;
rom[231] = 12'hccc;
rom[232] = 12'hccc;
rom[233] = 12'h007;
rom[234] = 12'h007;
rom[235] = 12'h007;
rom[236] = 12'hccc;
rom[237] = 12'hccc;
rom[238] = 12'hccc;
rom[239] = 12'hccc;
rom[240] = 12'hccc;
rom[241] = 12'hccc;
rom[242] = 12'hccc;
rom[243] = 12'hccc;
rom[244] = 12'hccc;
rom[245] = 12'hccc;
rom[246] = 12'hccc;
rom[247] = 12'hccc;
rom[248] = 12'hccc;
rom[249] = 12'h777;
rom[250] = 12'h777;
rom[251] = 12'hccc;
rom[252] = 12'hccc;
rom[253] = 12'hccc;
rom[254] = 12'hccc;
rom[255] = 12'hccc;
rom[256] = 12'hccc;
rom[257] = 12'hccc;
rom[258] = 12'h007;
rom[259] = 12'h007;
rom[260] = 12'h007;
rom[261] = 12'hccc;
rom[262] = 12'hccc;
rom[263] = 12'hccc;
rom[264] = 12'hccc;
rom[265] = 12'hccc;
rom[266] = 12'hccc;
rom[267] = 12'hccc;
rom[268] = 12'hccc;
rom[269] = 12'hccc;
rom[270] = 12'hccc;
rom[271] = 12'hccc;
rom[272] = 12'hccc;
rom[273] = 12'hccc;
rom[274] = 12'h777;
rom[275] = 12'h777;
rom[276] = 12'hccc;
rom[277] = 12'hccc;
rom[278] = 12'hccc;
rom[279] = 12'hccc;
rom[280] = 12'hccc;
rom[281] = 12'hccc;
rom[282] = 12'hccc;
rom[283] = 12'h007;
rom[284] = 12'h007;
rom[285] = 12'h007;
rom[286] = 12'h007;
rom[287] = 12'h007;
rom[288] = 12'h007;
rom[289] = 12'h007;
rom[290] = 12'h007;
rom[291] = 12'h007;
rom[292] = 12'hccc;
rom[293] = 12'hccc;
rom[294] = 12'hccc;
rom[295] = 12'hccc;
rom[296] = 12'hccc;
rom[297] = 12'hccc;
rom[298] = 12'hccc;
rom[299] = 12'h777;
rom[300] = 12'h777;
rom[301] = 12'hccc;
rom[302] = 12'hccc;
rom[303] = 12'hccc;
rom[304] = 12'hccc;
rom[305] = 12'hccc;
rom[306] = 12'hccc;
rom[307] = 12'hccc;
rom[308] = 12'h007;
rom[309] = 12'h007;
rom[310] = 12'h007;
rom[311] = 12'h007;
rom[312] = 12'h007;
rom[313] = 12'h007;
rom[314] = 12'h007;
rom[315] = 12'h007;
rom[316] = 12'h007;
rom[317] = 12'h007;
rom[318] = 12'hccc;
rom[319] = 12'hccc;
rom[320] = 12'hccc;
rom[321] = 12'hccc;
rom[322] = 12'hccc;
rom[323] = 12'hccc;
rom[324] = 12'h777;
rom[325] = 12'h777;
rom[326] = 12'hccc;
rom[327] = 12'hccc;
rom[328] = 12'hccc;
rom[329] = 12'hccc;
rom[330] = 12'hccc;
rom[331] = 12'hccc;
rom[332] = 12'hccc;
rom[333] = 12'hccc;
rom[334] = 12'hccc;
rom[335] = 12'hccc;
rom[336] = 12'hccc;
rom[337] = 12'hccc;
rom[338] = 12'hccc;
rom[339] = 12'hccc;
rom[340] = 12'h007;
rom[341] = 12'h007;
rom[342] = 12'h007;
rom[343] = 12'hccc;
rom[344] = 12'hccc;
rom[345] = 12'hccc;
rom[346] = 12'hccc;
rom[347] = 12'hccc;
rom[348] = 12'hccc;
rom[349] = 12'h777;
rom[350] = 12'h777;
rom[351] = 12'hccc;
rom[352] = 12'hccc;
rom[353] = 12'hccc;
rom[354] = 12'hccc;
rom[355] = 12'hccc;
rom[356] = 12'hccc;
rom[357] = 12'hccc;
rom[358] = 12'hccc;
rom[359] = 12'hccc;
rom[360] = 12'hccc;
rom[361] = 12'hccc;
rom[362] = 12'hccc;
rom[363] = 12'hccc;
rom[364] = 12'hccc;
rom[365] = 12'h007;
rom[366] = 12'h007;
rom[367] = 12'h007;
rom[368] = 12'hccc;
rom[369] = 12'hccc;
rom[370] = 12'hccc;
rom[371] = 12'hccc;
rom[372] = 12'hccc;
rom[373] = 12'hccc;
rom[374] = 12'h777;
rom[375] = 12'h777;
rom[376] = 12'hccc;
rom[377] = 12'hccc;
rom[378] = 12'hccc;
rom[379] = 12'hccc;
rom[380] = 12'hccc;
rom[381] = 12'hccc;
rom[382] = 12'hccc;
rom[383] = 12'h007;
rom[384] = 12'h007;
rom[385] = 12'h007;
rom[386] = 12'h007;
rom[387] = 12'h007;
rom[388] = 12'h007;
rom[389] = 12'h007;
rom[390] = 12'h007;
rom[391] = 12'h007;
rom[392] = 12'h007;
rom[393] = 12'hccc;
rom[394] = 12'hccc;
rom[395] = 12'hccc;
rom[396] = 12'hccc;
rom[397] = 12'hccc;
rom[398] = 12'hccc;
rom[399] = 12'h777;
rom[400] = 12'h777;
rom[401] = 12'hccc;
rom[402] = 12'hccc;
rom[403] = 12'hccc;
rom[404] = 12'hccc;
rom[405] = 12'hccc;
rom[406] = 12'hccc;
rom[407] = 12'hccc;
rom[408] = 12'h007;
rom[409] = 12'h007;
rom[410] = 12'h007;
rom[411] = 12'h007;
rom[412] = 12'h007;
rom[413] = 12'h007;
rom[414] = 12'h007;
rom[415] = 12'h007;
rom[416] = 12'h007;
rom[417] = 12'hccc;
rom[418] = 12'hccc;
rom[419] = 12'hccc;
rom[420] = 12'hccc;
rom[421] = 12'hccc;
rom[422] = 12'hccc;
rom[423] = 12'hccc;
rom[424] = 12'h777;
rom[425] = 12'h777;
rom[426] = 12'hccc;
rom[427] = 12'hccc;
rom[428] = 12'hccc;
rom[429] = 12'hccc;
rom[430] = 12'hccc;
rom[431] = 12'hccc;
rom[432] = 12'hccc;
rom[433] = 12'hccc;
rom[434] = 12'hccc;
rom[435] = 12'hccc;
rom[436] = 12'hccc;
rom[437] = 12'hccc;
rom[438] = 12'hccc;
rom[439] = 12'hccc;
rom[440] = 12'hbbb;
rom[441] = 12'hccc;
rom[442] = 12'hccc;
rom[443] = 12'hccc;
rom[444] = 12'hccc;
rom[445] = 12'hccc;
rom[446] = 12'hccc;
rom[447] = 12'hccc;
rom[448] = 12'hccc;
rom[449] = 12'h777;
rom[450] = 12'h777;
rom[451] = 12'hccc;
rom[452] = 12'hccc;
rom[453] = 12'hccc;
rom[454] = 12'hccc;
rom[455] = 12'hccc;
rom[456] = 12'hccc;
rom[457] = 12'hccc;
rom[458] = 12'hccc;
rom[459] = 12'hccc;
rom[460] = 12'hccc;
rom[461] = 12'hccc;
rom[462] = 12'hccc;
rom[463] = 12'hccc;
rom[464] = 12'hccc;
rom[465] = 12'hbbb;
rom[466] = 12'hccc;
rom[467] = 12'hccc;
rom[468] = 12'hccc;
rom[469] = 12'hccc;
rom[470] = 12'hccc;
rom[471] = 12'hccc;
rom[472] = 12'hccc;
rom[473] = 12'hccc;
rom[474] = 12'h777;
rom[475] = 12'h777;
rom[476] = 12'hccc;
rom[477] = 12'hccc;
rom[478] = 12'hccc;
rom[479] = 12'hccc;
rom[480] = 12'hccc;
rom[481] = 12'hccc;
rom[482] = 12'hccc;
rom[483] = 12'hccc;
rom[484] = 12'hccc;
rom[485] = 12'hccc;
rom[486] = 12'hccc;
rom[487] = 12'hccc;
rom[488] = 12'hccc;
rom[489] = 12'hccc;
rom[490] = 12'hccc;
rom[491] = 12'hccc;
rom[492] = 12'hccc;
rom[493] = 12'hccc;
rom[494] = 12'hccc;
rom[495] = 12'hccc;
rom[496] = 12'hccc;
rom[497] = 12'hccc;
rom[498] = 12'hccc;
rom[499] = 12'h777;
rom[500] = 12'h777;
rom[501] = 12'hccc;
rom[502] = 12'hccc;
rom[503] = 12'hccc;
rom[504] = 12'hccc;
rom[505] = 12'hccc;
rom[506] = 12'hccc;
rom[507] = 12'hccc;
rom[508] = 12'hccc;
rom[509] = 12'hccc;
rom[510] = 12'hccc;
rom[511] = 12'hccc;
rom[512] = 12'hccc;
rom[513] = 12'hccc;
rom[514] = 12'hccc;
rom[515] = 12'hccc;
rom[516] = 12'hccc;
rom[517] = 12'hccc;
rom[518] = 12'hccc;
rom[519] = 12'hccc;
rom[520] = 12'hccc;
rom[521] = 12'hccc;
rom[522] = 12'hccc;
rom[523] = 12'hccc;
rom[524] = 12'h777;
rom[525] = 12'h777;
rom[526] = 12'hccc;
rom[527] = 12'hccc;
rom[528] = 12'hccc;
rom[529] = 12'hccc;
rom[530] = 12'hccc;
rom[531] = 12'hccc;
rom[532] = 12'hccc;
rom[533] = 12'hccc;
rom[534] = 12'hccc;
rom[535] = 12'hccc;
rom[536] = 12'hccc;
rom[537] = 12'hccc;
rom[538] = 12'hccc;
rom[539] = 12'hccc;
rom[540] = 12'hccc;
rom[541] = 12'hccc;
rom[542] = 12'hccc;
rom[543] = 12'hccc;
rom[544] = 12'hccc;
rom[545] = 12'hccc;
rom[546] = 12'hccc;
rom[547] = 12'hccc;
rom[548] = 12'hccc;
rom[549] = 12'h777;
rom[550] = 12'h777;
rom[551] = 12'hccc;
rom[552] = 12'hccc;
rom[553] = 12'hccc;
rom[554] = 12'hccc;
rom[555] = 12'hccc;
rom[556] = 12'hccc;
rom[557] = 12'hccc;
rom[558] = 12'hccc;
rom[559] = 12'hccc;
rom[560] = 12'hccc;
rom[561] = 12'hccc;
rom[562] = 12'hccc;
rom[563] = 12'hccc;
rom[564] = 12'hccc;
rom[565] = 12'hccc;
rom[566] = 12'hccc;
rom[567] = 12'hccc;
rom[568] = 12'hccc;
rom[569] = 12'hccc;
rom[570] = 12'hccc;
rom[571] = 12'hccc;
rom[572] = 12'hccc;
rom[573] = 12'hccc;
rom[574] = 12'h777;
rom[575] = 12'h777;
rom[576] = 12'hccc;
rom[577] = 12'hccc;
rom[578] = 12'hccc;
rom[579] = 12'hccc;
rom[580] = 12'hccc;
rom[581] = 12'hccc;
rom[582] = 12'hccc;
rom[583] = 12'hccc;
rom[584] = 12'hccc;
rom[585] = 12'hccc;
rom[586] = 12'hccc;
rom[587] = 12'hccc;
rom[588] = 12'hccc;
rom[589] = 12'hccc;
rom[590] = 12'hccc;
rom[591] = 12'hccc;
rom[592] = 12'hccc;
rom[593] = 12'hccc;
rom[594] = 12'hccc;
rom[595] = 12'hccc;
rom[596] = 12'hccc;
rom[597] = 12'hccc;
rom[598] = 12'hccc;
rom[599] = 12'h777;
rom[600] = 12'h777;
rom[601] = 12'h777;
rom[602] = 12'h777;
rom[603] = 12'h777;
rom[604] = 12'h777;
rom[605] = 12'h777;
rom[606] = 12'h777;
rom[607] = 12'h777;
rom[608] = 12'h777;
rom[609] = 12'h777;
rom[610] = 12'h777;
rom[611] = 12'h777;
rom[612] = 12'h777;
rom[613] = 12'h777;
rom[614] = 12'h777;
rom[615] = 12'h777;
rom[616] = 12'h777;
rom[617] = 12'h777;
rom[618] = 12'h777;
rom[619] = 12'h777;
rom[620] = 12'h777;
rom[621] = 12'h777;
rom[622] = 12'h777;
rom[623] = 12'h777;
rom[624] = 12'h777;
  end
  endmodule

  module tile_six_rom (                       //клетка с шесёркой
  input  wire    [13:0]     addr,
  output wire    [11:0]     word
);

  logic [11:0] rom [(25 * 25)];

  assign word = rom[addr];

  initial begin
rom[0] = 12'h777;
rom[1] = 12'h777;
rom[2] = 12'h777;
rom[3] = 12'h777;
rom[4] = 12'h777;
rom[5] = 12'h777;
rom[6] = 12'h777;
rom[7] = 12'h777;
rom[8] = 12'h777;
rom[9] = 12'h777;
rom[10] = 12'h777;
rom[11] = 12'h777;
rom[12] = 12'h777;
rom[13] = 12'h777;
rom[14] = 12'h777;
rom[15] = 12'h777;
rom[16] = 12'h777;
rom[17] = 12'h777;
rom[18] = 12'h777;
rom[19] = 12'h777;
rom[20] = 12'h777;
rom[21] = 12'h777;
rom[22] = 12'h777;
rom[23] = 12'h777;
rom[24] = 12'h777;
rom[25] = 12'h777;
rom[26] = 12'hccc;
rom[27] = 12'hccc;
rom[28] = 12'hccc;
rom[29] = 12'hccc;
rom[30] = 12'hccc;
rom[31] = 12'hccc;
rom[32] = 12'hccc;
rom[33] = 12'hccc;
rom[34] = 12'hccc;
rom[35] = 12'hccc;
rom[36] = 12'hccc;
rom[37] = 12'hccc;
rom[38] = 12'hccc;
rom[39] = 12'hccc;
rom[40] = 12'hccc;
rom[41] = 12'hccc;
rom[42] = 12'hccc;
rom[43] = 12'hccc;
rom[44] = 12'hccc;
rom[45] = 12'hccc;
rom[46] = 12'hccc;
rom[47] = 12'hccc;
rom[48] = 12'hccc;
rom[49] = 12'h777;
rom[50] = 12'h777;
rom[51] = 12'hccc;
rom[52] = 12'hccc;
rom[53] = 12'hccc;
rom[54] = 12'hccc;
rom[55] = 12'hccc;
rom[56] = 12'hccc;
rom[57] = 12'hccc;
rom[58] = 12'hccc;
rom[59] = 12'hccc;
rom[60] = 12'hccc;
rom[61] = 12'hccc;
rom[62] = 12'hccc;
rom[63] = 12'hccc;
rom[64] = 12'hccc;
rom[65] = 12'hccc;
rom[66] = 12'hccc;
rom[67] = 12'hccc;
rom[68] = 12'hccc;
rom[69] = 12'hccc;
rom[70] = 12'hccc;
rom[71] = 12'hccc;
rom[72] = 12'hccc;
rom[73] = 12'hccc;
rom[74] = 12'h777;
rom[75] = 12'h777;
rom[76] = 12'hccc;
rom[77] = 12'hccc;
rom[78] = 12'hccc;
rom[79] = 12'hccc;
rom[80] = 12'hccc;
rom[81] = 12'hccc;
rom[82] = 12'hccc;
rom[83] = 12'hccc;
rom[84] = 12'hccc;
rom[85] = 12'hccc;
rom[86] = 12'hccc;
rom[87] = 12'hccc;
rom[88] = 12'hccc;
rom[89] = 12'hccc;
rom[90] = 12'hccc;
rom[91] = 12'hccc;
rom[92] = 12'hccc;
rom[93] = 12'hccc;
rom[94] = 12'hccc;
rom[95] = 12'hccc;
rom[96] = 12'hccc;
rom[97] = 12'hccc;
rom[98] = 12'hccc;
rom[99] = 12'h777;
rom[100] = 12'h777;
rom[101] = 12'hccc;
rom[102] = 12'hccc;
rom[103] = 12'hccc;
rom[104] = 12'hccc;
rom[105] = 12'hccc;
rom[106] = 12'hccc;
rom[107] = 12'hccc;
rom[108] = 12'hccc;
rom[109] = 12'hccc;
rom[110] = 12'hccc;
rom[111] = 12'hccc;
rom[112] = 12'hccc;
rom[113] = 12'hccc;
rom[114] = 12'hccc;
rom[115] = 12'hccc;
rom[116] = 12'hccc;
rom[117] = 12'hccc;
rom[118] = 12'hccc;
rom[119] = 12'hccc;
rom[120] = 12'hccc;
rom[121] = 12'hccc;
rom[122] = 12'hccc;
rom[123] = 12'hccc;
rom[124] = 12'h777;
rom[125] = 12'h777;
rom[126] = 12'hccc;
rom[127] = 12'hccc;
rom[128] = 12'hccc;
rom[129] = 12'hccc;
rom[130] = 12'hccc;
rom[131] = 12'hccc;
rom[132] = 12'hccc;
rom[133] = 12'hccc;
rom[134] = 12'hccc;
rom[135] = 12'hccc;
rom[136] = 12'hccc;
rom[137] = 12'hccc;
rom[138] = 12'hccc;
rom[139] = 12'hccc;
rom[140] = 12'hccc;
rom[141] = 12'hccc;
rom[142] = 12'hccc;
rom[143] = 12'hccc;
rom[144] = 12'hccc;
rom[145] = 12'hccc;
rom[146] = 12'hccc;
rom[147] = 12'hccc;
rom[148] = 12'hccc;
rom[149] = 12'h777;
rom[150] = 12'h777;
rom[151] = 12'hccc;
rom[152] = 12'hccc;
rom[153] = 12'hccc;
rom[154] = 12'hccc;
rom[155] = 12'hccc;
rom[156] = 12'hccc;
rom[157] = 12'hccc;
rom[158] = 12'hccc;
rom[159] = 12'hccc;
rom[160] = 12'hccc;
rom[161] = 12'hccc;
rom[162] = 12'hccc;
rom[163] = 12'hccc;
rom[164] = 12'hccc;
rom[165] = 12'hccc;
rom[166] = 12'hccc;
rom[167] = 12'hccc;
rom[168] = 12'hccc;
rom[169] = 12'hccc;
rom[170] = 12'hccc;
rom[171] = 12'hccc;
rom[172] = 12'hccc;
rom[173] = 12'hccc;
rom[174] = 12'h777;
rom[175] = 12'h777;
rom[176] = 12'hccc;
rom[177] = 12'hccc;
rom[178] = 12'hccc;
rom[179] = 12'hccc;
rom[180] = 12'hccc;
rom[181] = 12'hccc;
rom[182] = 12'hccc;
rom[183] = 12'hccc;
rom[184] = 12'h770;
rom[185] = 12'h770;
rom[186] = 12'h770;
rom[187] = 12'h770;
rom[188] = 12'h770;
rom[189] = 12'h770;
rom[190] = 12'h770;
rom[191] = 12'h770;
rom[192] = 12'hccc;
rom[193] = 12'hccc;
rom[194] = 12'hccc;
rom[195] = 12'hccc;
rom[196] = 12'hccc;
rom[197] = 12'hccc;
rom[198] = 12'hccc;
rom[199] = 12'h777;
rom[200] = 12'h777;
rom[201] = 12'hccc;
rom[202] = 12'hccc;
rom[203] = 12'hccc;
rom[204] = 12'hccc;
rom[205] = 12'hccc;
rom[206] = 12'hccc;
rom[207] = 12'hccc;
rom[208] = 12'h770;
rom[209] = 12'h770;
rom[210] = 12'h770;
rom[211] = 12'h770;
rom[212] = 12'h770;
rom[213] = 12'h770;
rom[214] = 12'h770;
rom[215] = 12'h770;
rom[216] = 12'h770;
rom[217] = 12'hccc;
rom[218] = 12'hccc;
rom[219] = 12'hccc;
rom[220] = 12'hccc;
rom[221] = 12'hccc;
rom[222] = 12'hccc;
rom[223] = 12'hccc;
rom[224] = 12'h777;
rom[225] = 12'h777;
rom[226] = 12'hccc;
rom[227] = 12'hccc;
rom[228] = 12'hccc;
rom[229] = 12'hccc;
rom[230] = 12'hccc;
rom[231] = 12'hccc;
rom[232] = 12'hccc;
rom[233] = 12'h770;
rom[234] = 12'h770;
rom[235] = 12'h770;
rom[236] = 12'hccc;
rom[237] = 12'hccc;
rom[238] = 12'hccc;
rom[239] = 12'hccc;
rom[240] = 12'hccc;
rom[241] = 12'hccc;
rom[242] = 12'hccc;
rom[243] = 12'hccc;
rom[244] = 12'hccc;
rom[245] = 12'hccc;
rom[246] = 12'hccc;
rom[247] = 12'hccc;
rom[248] = 12'hccc;
rom[249] = 12'h777;
rom[250] = 12'h777;
rom[251] = 12'hccc;
rom[252] = 12'hccc;
rom[253] = 12'hccc;
rom[254] = 12'hccc;
rom[255] = 12'hccc;
rom[256] = 12'hccc;
rom[257] = 12'hccc;
rom[258] = 12'h770;
rom[259] = 12'h770;
rom[260] = 12'h770;
rom[261] = 12'hccc;
rom[262] = 12'hccc;
rom[263] = 12'hccc;
rom[264] = 12'hccc;
rom[265] = 12'hccc;
rom[266] = 12'hccc;
rom[267] = 12'hccc;
rom[268] = 12'hccc;
rom[269] = 12'hccc;
rom[270] = 12'hccc;
rom[271] = 12'hccc;
rom[272] = 12'hccc;
rom[273] = 12'hccc;
rom[274] = 12'h777;
rom[275] = 12'h777;
rom[276] = 12'hccc;
rom[277] = 12'hccc;
rom[278] = 12'hccc;
rom[279] = 12'hccc;
rom[280] = 12'hccc;
rom[281] = 12'hccc;
rom[282] = 12'hccc;
rom[283] = 12'h770;
rom[284] = 12'h770;
rom[285] = 12'h770;
rom[286] = 12'h770;
rom[287] = 12'h770;
rom[288] = 12'h770;
rom[289] = 12'h770;
rom[290] = 12'h770;
rom[291] = 12'h770;
rom[292] = 12'hccc;
rom[293] = 12'hccc;
rom[294] = 12'hccc;
rom[295] = 12'hccc;
rom[296] = 12'hccc;
rom[297] = 12'hccc;
rom[298] = 12'hccc;
rom[299] = 12'h777;
rom[300] = 12'h777;
rom[301] = 12'hccc;
rom[302] = 12'hccc;
rom[303] = 12'hccc;
rom[304] = 12'hccc;
rom[305] = 12'hccc;
rom[306] = 12'hccc;
rom[307] = 12'hccc;
rom[308] = 12'h770;
rom[309] = 12'h770;
rom[310] = 12'h770;
rom[311] = 12'h770;
rom[312] = 12'h770;
rom[313] = 12'h770;
rom[314] = 12'h770;
rom[315] = 12'h770;
rom[316] = 12'h770;
rom[317] = 12'h770;
rom[318] = 12'hccc;
rom[319] = 12'hccc;
rom[320] = 12'hccc;
rom[321] = 12'hccc;
rom[322] = 12'hccc;
rom[323] = 12'hccc;
rom[324] = 12'h777;
rom[325] = 12'h777;
rom[326] = 12'hccc;
rom[327] = 12'hccc;
rom[328] = 12'hccc;
rom[329] = 12'hccc;
rom[330] = 12'hccc;
rom[331] = 12'hccc;
rom[332] = 12'hccc;
rom[333] = 12'h770;
rom[334] = 12'h770;
rom[335] = 12'h770;
rom[336] = 12'hccc;
rom[337] = 12'hccc;
rom[338] = 12'hccc;
rom[339] = 12'hccc;
rom[340] = 12'h770;
rom[341] = 12'h770;
rom[342] = 12'h770;
rom[343] = 12'hccc;
rom[344] = 12'hccc;
rom[345] = 12'hccc;
rom[346] = 12'hccc;
rom[347] = 12'hccc;
rom[348] = 12'hccc;
rom[349] = 12'h777;
rom[350] = 12'h777;
rom[351] = 12'hccc;
rom[352] = 12'hccc;
rom[353] = 12'hccc;
rom[354] = 12'hccc;
rom[355] = 12'hccc;
rom[356] = 12'hccc;
rom[357] = 12'hccc;
rom[358] = 12'h770;
rom[359] = 12'h770;
rom[360] = 12'h770;
rom[361] = 12'hccc;
rom[362] = 12'hccc;
rom[363] = 12'hccc;
rom[364] = 12'hccc;
rom[365] = 12'h770;
rom[366] = 12'h770;
rom[367] = 12'h770;
rom[368] = 12'hccc;
rom[369] = 12'hccc;
rom[370] = 12'hccc;
rom[371] = 12'hccc;
rom[372] = 12'hccc;
rom[373] = 12'hccc;
rom[374] = 12'h777;
rom[375] = 12'h777;
rom[376] = 12'hccc;
rom[377] = 12'hccc;
rom[378] = 12'hccc;
rom[379] = 12'hccc;
rom[380] = 12'hccc;
rom[381] = 12'hccc;
rom[382] = 12'hccc;
rom[383] = 12'h770;
rom[384] = 12'h770;
rom[385] = 12'h770;
rom[386] = 12'h770;
rom[387] = 12'h770;
rom[388] = 12'h770;
rom[389] = 12'h770;
rom[390] = 12'h770;
rom[391] = 12'h770;
rom[392] = 12'h770;
rom[393] = 12'hccc;
rom[394] = 12'hccc;
rom[395] = 12'hccc;
rom[396] = 12'hccc;
rom[397] = 12'hccc;
rom[398] = 12'hccc;
rom[399] = 12'h777;
rom[400] = 12'h777;
rom[401] = 12'hccc;
rom[402] = 12'hccc;
rom[403] = 12'hccc;
rom[404] = 12'hccc;
rom[405] = 12'hccc;
rom[406] = 12'hccc;
rom[407] = 12'hccc;
rom[408] = 12'hccc;
rom[409] = 12'h770;
rom[410] = 12'h770;
rom[411] = 12'h770;
rom[412] = 12'h770;
rom[413] = 12'h770;
rom[414] = 12'h770;
rom[415] = 12'h770;
rom[416] = 12'h770;
rom[417] = 12'hccc;
rom[418] = 12'hccc;
rom[419] = 12'hccc;
rom[420] = 12'hccc;
rom[421] = 12'hccc;
rom[422] = 12'hccc;
rom[423] = 12'hccc;
rom[424] = 12'h777;
rom[425] = 12'h777;
rom[426] = 12'hccc;
rom[427] = 12'hccc;
rom[428] = 12'hccc;
rom[429] = 12'hccc;
rom[430] = 12'hccc;
rom[431] = 12'hccc;
rom[432] = 12'hccc;
rom[433] = 12'hccc;
rom[434] = 12'hccc;
rom[435] = 12'hccc;
rom[436] = 12'hccc;
rom[437] = 12'hccc;
rom[438] = 12'hccc;
rom[439] = 12'hccc;
rom[440] = 12'hbbb;
rom[441] = 12'hccc;
rom[442] = 12'hccc;
rom[443] = 12'hccc;
rom[444] = 12'hccc;
rom[445] = 12'hccc;
rom[446] = 12'hccc;
rom[447] = 12'hccc;
rom[448] = 12'hccc;
rom[449] = 12'h777;
rom[450] = 12'h777;
rom[451] = 12'hccc;
rom[452] = 12'hccc;
rom[453] = 12'hccc;
rom[454] = 12'hccc;
rom[455] = 12'hccc;
rom[456] = 12'hccc;
rom[457] = 12'hccc;
rom[458] = 12'hccc;
rom[459] = 12'hccc;
rom[460] = 12'hccc;
rom[461] = 12'hccc;
rom[462] = 12'hccc;
rom[463] = 12'hccc;
rom[464] = 12'hccc;
rom[465] = 12'hbbb;
rom[466] = 12'hccc;
rom[467] = 12'hccc;
rom[468] = 12'hccc;
rom[469] = 12'hccc;
rom[470] = 12'hccc;
rom[471] = 12'hccc;
rom[472] = 12'hccc;
rom[473] = 12'hccc;
rom[474] = 12'h777;
rom[475] = 12'h777;
rom[476] = 12'hccc;
rom[477] = 12'hccc;
rom[478] = 12'hccc;
rom[479] = 12'hccc;
rom[480] = 12'hccc;
rom[481] = 12'hccc;
rom[482] = 12'hccc;
rom[483] = 12'hccc;
rom[484] = 12'hccc;
rom[485] = 12'hccc;
rom[486] = 12'hccc;
rom[487] = 12'hccc;
rom[488] = 12'hccc;
rom[489] = 12'hccc;
rom[490] = 12'hccc;
rom[491] = 12'hccc;
rom[492] = 12'hccc;
rom[493] = 12'hccc;
rom[494] = 12'hccc;
rom[495] = 12'hccc;
rom[496] = 12'hccc;
rom[497] = 12'hccc;
rom[498] = 12'hccc;
rom[499] = 12'h777;
rom[500] = 12'h777;
rom[501] = 12'hccc;
rom[502] = 12'hccc;
rom[503] = 12'hccc;
rom[504] = 12'hccc;
rom[505] = 12'hccc;
rom[506] = 12'hccc;
rom[507] = 12'hccc;
rom[508] = 12'hccc;
rom[509] = 12'hccc;
rom[510] = 12'hccc;
rom[511] = 12'hccc;
rom[512] = 12'hccc;
rom[513] = 12'hccc;
rom[514] = 12'hccc;
rom[515] = 12'hccc;
rom[516] = 12'hccc;
rom[517] = 12'hccc;
rom[518] = 12'hccc;
rom[519] = 12'hccc;
rom[520] = 12'hccc;
rom[521] = 12'hccc;
rom[522] = 12'hccc;
rom[523] = 12'hccc;
rom[524] = 12'h777;
rom[525] = 12'h777;
rom[526] = 12'hccc;
rom[527] = 12'hccc;
rom[528] = 12'hccc;
rom[529] = 12'hccc;
rom[530] = 12'hccc;
rom[531] = 12'hccc;
rom[532] = 12'hccc;
rom[533] = 12'hccc;
rom[534] = 12'hccc;
rom[535] = 12'hccc;
rom[536] = 12'hccc;
rom[537] = 12'hccc;
rom[538] = 12'hccc;
rom[539] = 12'hccc;
rom[540] = 12'hccc;
rom[541] = 12'hccc;
rom[542] = 12'hccc;
rom[543] = 12'hccc;
rom[544] = 12'hccc;
rom[545] = 12'hccc;
rom[546] = 12'hccc;
rom[547] = 12'hccc;
rom[548] = 12'hccc;
rom[549] = 12'h777;
rom[550] = 12'h777;
rom[551] = 12'hccc;
rom[552] = 12'hccc;
rom[553] = 12'hccc;
rom[554] = 12'hccc;
rom[555] = 12'hccc;
rom[556] = 12'hccc;
rom[557] = 12'hccc;
rom[558] = 12'hccc;
rom[559] = 12'hccc;
rom[560] = 12'hccc;
rom[561] = 12'hccc;
rom[562] = 12'hccc;
rom[563] = 12'hccc;
rom[564] = 12'hccc;
rom[565] = 12'hccc;
rom[566] = 12'hccc;
rom[567] = 12'hccc;
rom[568] = 12'hccc;
rom[569] = 12'hccc;
rom[570] = 12'hccc;
rom[571] = 12'hccc;
rom[572] = 12'hccc;
rom[573] = 12'hccc;
rom[574] = 12'h777;
rom[575] = 12'h777;
rom[576] = 12'hccc;
rom[577] = 12'hccc;
rom[578] = 12'hccc;
rom[579] = 12'hccc;
rom[580] = 12'hccc;
rom[581] = 12'hccc;
rom[582] = 12'hccc;
rom[583] = 12'hccc;
rom[584] = 12'hccc;
rom[585] = 12'hccc;
rom[586] = 12'hccc;
rom[587] = 12'hccc;
rom[588] = 12'hccc;
rom[589] = 12'hccc;
rom[590] = 12'hccc;
rom[591] = 12'hccc;
rom[592] = 12'hccc;
rom[593] = 12'hccc;
rom[594] = 12'hccc;
rom[595] = 12'hccc;
rom[596] = 12'hccc;
rom[597] = 12'hccc;
rom[598] = 12'hccc;
rom[599] = 12'h777;
rom[600] = 12'h777;
rom[601] = 12'h777;
rom[602] = 12'h777;
rom[603] = 12'h777;
rom[604] = 12'h777;
rom[605] = 12'h777;
rom[606] = 12'h777;
rom[607] = 12'h777;
rom[608] = 12'h777;
rom[609] = 12'h777;
rom[610] = 12'h777;
rom[611] = 12'h777;
rom[612] = 12'h777;
rom[613] = 12'h777;
rom[614] = 12'h777;
rom[615] = 12'h777;
rom[616] = 12'h777;
rom[617] = 12'h777;
rom[618] = 12'h777;
rom[619] = 12'h777;
rom[620] = 12'h777;
rom[621] = 12'h777;
rom[622] = 12'h777;
rom[623] = 12'h777;
rom[624] = 12'h777;
  end
  endmodule

  module tile_seven_rom (                       //клетка с семёркой
  input  wire    [13:0]     addr,
  output wire    [11:0]     word
);

  logic [11:0] rom [(25 * 25)];

  assign word = rom[addr];

  initial begin
rom[0] = 12'h777;
rom[1] = 12'h777;
rom[2] = 12'h777;
rom[3] = 12'h777;
rom[4] = 12'h777;
rom[5] = 12'h777;
rom[6] = 12'h777;
rom[7] = 12'h777;
rom[8] = 12'h777;
rom[9] = 12'h777;
rom[10] = 12'h777;
rom[11] = 12'h777;
rom[12] = 12'h777;
rom[13] = 12'h777;
rom[14] = 12'h777;
rom[15] = 12'h777;
rom[16] = 12'h777;
rom[17] = 12'h777;
rom[18] = 12'h777;
rom[19] = 12'h777;
rom[20] = 12'h777;
rom[21] = 12'h777;
rom[22] = 12'h777;
rom[23] = 12'h777;
rom[24] = 12'h777;
rom[25] = 12'h777;
rom[26] = 12'hccc;
rom[27] = 12'hccc;
rom[28] = 12'hccc;
rom[29] = 12'hccc;
rom[30] = 12'hccc;
rom[31] = 12'hccc;
rom[32] = 12'hccc;
rom[33] = 12'hccc;
rom[34] = 12'hccc;
rom[35] = 12'hccc;
rom[36] = 12'hccc;
rom[37] = 12'hccc;
rom[38] = 12'hccc;
rom[39] = 12'hccc;
rom[40] = 12'hccc;
rom[41] = 12'hccc;
rom[42] = 12'hccc;
rom[43] = 12'hccc;
rom[44] = 12'hccc;
rom[45] = 12'hccc;
rom[46] = 12'hccc;
rom[47] = 12'hccc;
rom[48] = 12'hccc;
rom[49] = 12'h777;
rom[50] = 12'h777;
rom[51] = 12'hccc;
rom[52] = 12'hccc;
rom[53] = 12'hccc;
rom[54] = 12'hccc;
rom[55] = 12'hccc;
rom[56] = 12'hccc;
rom[57] = 12'hccc;
rom[58] = 12'hccc;
rom[59] = 12'hccc;
rom[60] = 12'hccc;
rom[61] = 12'hccc;
rom[62] = 12'hccc;
rom[63] = 12'hccc;
rom[64] = 12'hccc;
rom[65] = 12'hccc;
rom[66] = 12'hccc;
rom[67] = 12'hccc;
rom[68] = 12'hccc;
rom[69] = 12'hccc;
rom[70] = 12'hccc;
rom[71] = 12'hccc;
rom[72] = 12'hccc;
rom[73] = 12'hccc;
rom[74] = 12'h777;
rom[75] = 12'h777;
rom[76] = 12'hccc;
rom[77] = 12'hccc;
rom[78] = 12'hccc;
rom[79] = 12'hccc;
rom[80] = 12'hccc;
rom[81] = 12'hccc;
rom[82] = 12'hccc;
rom[83] = 12'hccc;
rom[84] = 12'hccc;
rom[85] = 12'hccc;
rom[86] = 12'hccc;
rom[87] = 12'hccc;
rom[88] = 12'hccc;
rom[89] = 12'hccc;
rom[90] = 12'hccc;
rom[91] = 12'hccc;
rom[92] = 12'hccc;
rom[93] = 12'hccc;
rom[94] = 12'hccc;
rom[95] = 12'hccc;
rom[96] = 12'hccc;
rom[97] = 12'hccc;
rom[98] = 12'hccc;
rom[99] = 12'h777;
rom[100] = 12'h777;
rom[101] = 12'hccc;
rom[102] = 12'hccc;
rom[103] = 12'hccc;
rom[104] = 12'hccc;
rom[105] = 12'hccc;
rom[106] = 12'hccc;
rom[107] = 12'hccc;
rom[108] = 12'hccc;
rom[109] = 12'hccc;
rom[110] = 12'hccc;
rom[111] = 12'hccc;
rom[112] = 12'hccc;
rom[113] = 12'hccc;
rom[114] = 12'hccc;
rom[115] = 12'hccc;
rom[116] = 12'hccc;
rom[117] = 12'hccc;
rom[118] = 12'hccc;
rom[119] = 12'hccc;
rom[120] = 12'hccc;
rom[121] = 12'hccc;
rom[122] = 12'hccc;
rom[123] = 12'hccc;
rom[124] = 12'h777;
rom[125] = 12'h777;
rom[126] = 12'hccc;
rom[127] = 12'hccc;
rom[128] = 12'hccc;
rom[129] = 12'hccc;
rom[130] = 12'hccc;
rom[131] = 12'hccc;
rom[132] = 12'hccc;
rom[133] = 12'hccc;
rom[134] = 12'hccc;
rom[135] = 12'hccc;
rom[136] = 12'hccc;
rom[137] = 12'hccc;
rom[138] = 12'hccc;
rom[139] = 12'hccc;
rom[140] = 12'hccc;
rom[141] = 12'hccc;
rom[142] = 12'hccc;
rom[143] = 12'hccc;
rom[144] = 12'hccc;
rom[145] = 12'hccc;
rom[146] = 12'hccc;
rom[147] = 12'hccc;
rom[148] = 12'hccc;
rom[149] = 12'h777;
rom[150] = 12'h777;
rom[151] = 12'hccc;
rom[152] = 12'hccc;
rom[153] = 12'hccc;
rom[154] = 12'hccc;
rom[155] = 12'hccc;
rom[156] = 12'hccc;
rom[157] = 12'hccc;
rom[158] = 12'hccc;
rom[159] = 12'hccc;
rom[160] = 12'hccc;
rom[161] = 12'hccc;
rom[162] = 12'hccc;
rom[163] = 12'hccc;
rom[164] = 12'hccc;
rom[165] = 12'hccc;
rom[166] = 12'hccc;
rom[167] = 12'hccc;
rom[168] = 12'hccc;
rom[169] = 12'hccc;
rom[170] = 12'hccc;
rom[171] = 12'hccc;
rom[172] = 12'hccc;
rom[173] = 12'hccc;
rom[174] = 12'h777;
rom[175] = 12'h777;
rom[176] = 12'hccc;
rom[177] = 12'hccc;
rom[178] = 12'hccc;
rom[179] = 12'hccc;
rom[180] = 12'hccc;
rom[181] = 12'hccc;
rom[182] = 12'hccc;
rom[183] = 12'h000;
rom[184] = 12'h000;
rom[185] = 12'h000;
rom[186] = 12'h000;
rom[187] = 12'h000;
rom[188] = 12'h000;
rom[189] = 12'h000;
rom[190] = 12'h000;
rom[191] = 12'h000;
rom[192] = 12'h000;
rom[193] = 12'hccc;
rom[194] = 12'hccc;
rom[195] = 12'hccc;
rom[196] = 12'hccc;
rom[197] = 12'hccc;
rom[198] = 12'hccc;
rom[199] = 12'h777;
rom[200] = 12'h777;
rom[201] = 12'hccc;
rom[202] = 12'hccc;
rom[203] = 12'hccc;
rom[204] = 12'hccc;
rom[205] = 12'hccc;
rom[206] = 12'hccc;
rom[207] = 12'hccc;
rom[208] = 12'h000;
rom[209] = 12'h000;
rom[210] = 12'h000;
rom[211] = 12'h000;
rom[212] = 12'h000;
rom[213] = 12'h000;
rom[214] = 12'h000;
rom[215] = 12'h000;
rom[216] = 12'h000;
rom[217] = 12'h000;
rom[218] = 12'hccc;
rom[219] = 12'hccc;
rom[220] = 12'hccc;
rom[221] = 12'hccc;
rom[222] = 12'hccc;
rom[223] = 12'hccc;
rom[224] = 12'h777;
rom[225] = 12'h777;
rom[226] = 12'hccc;
rom[227] = 12'hccc;
rom[228] = 12'hccc;
rom[229] = 12'hccc;
rom[230] = 12'hccc;
rom[231] = 12'hccc;
rom[232] = 12'hccc;
rom[233] = 12'hccc;
rom[234] = 12'hccc;
rom[235] = 12'hccc;
rom[236] = 12'hccc;
rom[237] = 12'hccc;
rom[238] = 12'hccc;
rom[239] = 12'hccc;
rom[240] = 12'h000;
rom[241] = 12'h000;
rom[242] = 12'h000;
rom[243] = 12'hccc;
rom[244] = 12'hccc;
rom[245] = 12'hccc;
rom[246] = 12'hccc;
rom[247] = 12'hccc;
rom[248] = 12'hccc;
rom[249] = 12'h777;
rom[250] = 12'h777;
rom[251] = 12'hccc;
rom[252] = 12'hccc;
rom[253] = 12'hccc;
rom[254] = 12'hccc;
rom[255] = 12'hccc;
rom[256] = 12'hccc;
rom[257] = 12'hccc;
rom[258] = 12'hccc;
rom[259] = 12'hccc;
rom[260] = 12'hccc;
rom[261] = 12'hccc;
rom[262] = 12'hccc;
rom[263] = 12'hccc;
rom[264] = 12'hccc;
rom[265] = 12'h000;
rom[266] = 12'h000;
rom[267] = 12'h000;
rom[268] = 12'hccc;
rom[269] = 12'hccc;
rom[270] = 12'hccc;
rom[271] = 12'hccc;
rom[272] = 12'hccc;
rom[273] = 12'hccc;
rom[274] = 12'h777;
rom[275] = 12'h777;
rom[276] = 12'hccc;
rom[277] = 12'hccc;
rom[278] = 12'hccc;
rom[279] = 12'hccc;
rom[280] = 12'hccc;
rom[281] = 12'hccc;
rom[282] = 12'hccc;
rom[283] = 12'hccc;
rom[284] = 12'hccc;
rom[285] = 12'hccc;
rom[286] = 12'hccc;
rom[287] = 12'hccc;
rom[288] = 12'hccc;
rom[289] = 12'h000;
rom[290] = 12'h000;
rom[291] = 12'h000;
rom[292] = 12'hccc;
rom[293] = 12'hccc;
rom[294] = 12'hccc;
rom[295] = 12'hccc;
rom[296] = 12'hccc;
rom[297] = 12'hccc;
rom[298] = 12'hccc;
rom[299] = 12'h777;
rom[300] = 12'h777;
rom[301] = 12'hccc;
rom[302] = 12'hccc;
rom[303] = 12'hccc;
rom[304] = 12'hccc;
rom[305] = 12'hccc;
rom[306] = 12'hccc;
rom[307] = 12'hccc;
rom[308] = 12'hccc;
rom[309] = 12'hccc;
rom[310] = 12'hccc;
rom[311] = 12'hccc;
rom[312] = 12'hccc;
rom[313] = 12'hccc;
rom[314] = 12'h000;
rom[315] = 12'h000;
rom[316] = 12'h000;
rom[317] = 12'hccc;
rom[318] = 12'hccc;
rom[319] = 12'hccc;
rom[320] = 12'hccc;
rom[321] = 12'hccc;
rom[322] = 12'hccc;
rom[323] = 12'hccc;
rom[324] = 12'h777;
rom[325] = 12'h777;
rom[326] = 12'hccc;
rom[327] = 12'hccc;
rom[328] = 12'hccc;
rom[329] = 12'hccc;
rom[330] = 12'hccc;
rom[331] = 12'hccc;
rom[332] = 12'hccc;
rom[333] = 12'hccc;
rom[334] = 12'hccc;
rom[335] = 12'hccc;
rom[336] = 12'hccc;
rom[337] = 12'hccc;
rom[338] = 12'h000;
rom[339] = 12'h000;
rom[340] = 12'h000;
rom[341] = 12'hccc;
rom[342] = 12'hccc;
rom[343] = 12'hccc;
rom[344] = 12'hccc;
rom[345] = 12'hccc;
rom[346] = 12'hccc;
rom[347] = 12'hccc;
rom[348] = 12'hccc;
rom[349] = 12'h777;
rom[350] = 12'h777;
rom[351] = 12'hccc;
rom[352] = 12'hccc;
rom[353] = 12'hccc;
rom[354] = 12'hccc;
rom[355] = 12'hccc;
rom[356] = 12'hccc;
rom[357] = 12'hccc;
rom[358] = 12'hccc;
rom[359] = 12'hccc;
rom[360] = 12'hccc;
rom[361] = 12'hccc;
rom[362] = 12'hccc;
rom[363] = 12'h000;
rom[364] = 12'h000;
rom[365] = 12'h000;
rom[366] = 12'hccc;
rom[367] = 12'hccc;
rom[368] = 12'hccc;
rom[369] = 12'hccc;
rom[370] = 12'hccc;
rom[371] = 12'hccc;
rom[372] = 12'hccc;
rom[373] = 12'hccc;
rom[374] = 12'h777;
rom[375] = 12'h777;
rom[376] = 12'hccc;
rom[377] = 12'hccc;
rom[378] = 12'hccc;
rom[379] = 12'hccc;
rom[380] = 12'hccc;
rom[381] = 12'hccc;
rom[382] = 12'hccc;
rom[383] = 12'hccc;
rom[384] = 12'hccc;
rom[385] = 12'hccc;
rom[386] = 12'hccc;
rom[387] = 12'h000;
rom[388] = 12'h000;
rom[389] = 12'h000;
rom[390] = 12'hccc;
rom[391] = 12'hccc;
rom[392] = 12'hccc;
rom[393] = 12'hccc;
rom[394] = 12'hccc;
rom[395] = 12'hccc;
rom[396] = 12'hccc;
rom[397] = 12'hccc;
rom[398] = 12'hccc;
rom[399] = 12'h777;
rom[400] = 12'h777;
rom[401] = 12'hccc;
rom[402] = 12'hccc;
rom[403] = 12'hccc;
rom[404] = 12'hccc;
rom[405] = 12'hccc;
rom[406] = 12'hccc;
rom[407] = 12'hccc;
rom[408] = 12'hccc;
rom[409] = 12'hccc;
rom[410] = 12'hccc;
rom[411] = 12'hccc;
rom[412] = 12'h000;
rom[413] = 12'h000;
rom[414] = 12'h000;
rom[415] = 12'hccc;
rom[416] = 12'hccc;
rom[417] = 12'hccc;
rom[418] = 12'hccc;
rom[419] = 12'hccc;
rom[420] = 12'hccc;
rom[421] = 12'hccc;
rom[422] = 12'hccc;
rom[423] = 12'hccc;
rom[424] = 12'h777;
rom[425] = 12'h777;
rom[426] = 12'hccc;
rom[427] = 12'hccc;
rom[428] = 12'hccc;
rom[429] = 12'hccc;
rom[430] = 12'hccc;
rom[431] = 12'hccc;
rom[432] = 12'hccc;
rom[433] = 12'hccc;
rom[434] = 12'hccc;
rom[435] = 12'hccc;
rom[436] = 12'hccc;
rom[437] = 12'hccc;
rom[438] = 12'hccc;
rom[439] = 12'hccc;
rom[440] = 12'hbbb;
rom[441] = 12'hccc;
rom[442] = 12'hccc;
rom[443] = 12'hccc;
rom[444] = 12'hccc;
rom[445] = 12'hccc;
rom[446] = 12'hccc;
rom[447] = 12'hccc;
rom[448] = 12'hccc;
rom[449] = 12'h777;
rom[450] = 12'h777;
rom[451] = 12'hccc;
rom[452] = 12'hccc;
rom[453] = 12'hccc;
rom[454] = 12'hccc;
rom[455] = 12'hccc;
rom[456] = 12'hccc;
rom[457] = 12'hccc;
rom[458] = 12'hccc;
rom[459] = 12'hccc;
rom[460] = 12'hccc;
rom[461] = 12'hccc;
rom[462] = 12'hccc;
rom[463] = 12'hccc;
rom[464] = 12'hccc;
rom[465] = 12'hbbb;
rom[466] = 12'hccc;
rom[467] = 12'hccc;
rom[468] = 12'hccc;
rom[469] = 12'hccc;
rom[470] = 12'hccc;
rom[471] = 12'hccc;
rom[472] = 12'hccc;
rom[473] = 12'hccc;
rom[474] = 12'h777;
rom[475] = 12'h777;
rom[476] = 12'hccc;
rom[477] = 12'hccc;
rom[478] = 12'hccc;
rom[479] = 12'hccc;
rom[480] = 12'hccc;
rom[481] = 12'hccc;
rom[482] = 12'hccc;
rom[483] = 12'hccc;
rom[484] = 12'hccc;
rom[485] = 12'hccc;
rom[486] = 12'hccc;
rom[487] = 12'hccc;
rom[488] = 12'hccc;
rom[489] = 12'hccc;
rom[490] = 12'hccc;
rom[491] = 12'hccc;
rom[492] = 12'hccc;
rom[493] = 12'hccc;
rom[494] = 12'hccc;
rom[495] = 12'hccc;
rom[496] = 12'hccc;
rom[497] = 12'hccc;
rom[498] = 12'hccc;
rom[499] = 12'h777;
rom[500] = 12'h777;
rom[501] = 12'hccc;
rom[502] = 12'hccc;
rom[503] = 12'hccc;
rom[504] = 12'hccc;
rom[505] = 12'hccc;
rom[506] = 12'hccc;
rom[507] = 12'hccc;
rom[508] = 12'hccc;
rom[509] = 12'hccc;
rom[510] = 12'hccc;
rom[511] = 12'hccc;
rom[512] = 12'hccc;
rom[513] = 12'hccc;
rom[514] = 12'hccc;
rom[515] = 12'hccc;
rom[516] = 12'hccc;
rom[517] = 12'hccc;
rom[518] = 12'hccc;
rom[519] = 12'hccc;
rom[520] = 12'hccc;
rom[521] = 12'hccc;
rom[522] = 12'hccc;
rom[523] = 12'hccc;
rom[524] = 12'h777;
rom[525] = 12'h777;
rom[526] = 12'hccc;
rom[527] = 12'hccc;
rom[528] = 12'hccc;
rom[529] = 12'hccc;
rom[530] = 12'hccc;
rom[531] = 12'hccc;
rom[532] = 12'hccc;
rom[533] = 12'hccc;
rom[534] = 12'hccc;
rom[535] = 12'hccc;
rom[536] = 12'hccc;
rom[537] = 12'hccc;
rom[538] = 12'hccc;
rom[539] = 12'hccc;
rom[540] = 12'hccc;
rom[541] = 12'hccc;
rom[542] = 12'hccc;
rom[543] = 12'hccc;
rom[544] = 12'hccc;
rom[545] = 12'hccc;
rom[546] = 12'hccc;
rom[547] = 12'hccc;
rom[548] = 12'hccc;
rom[549] = 12'h777;
rom[550] = 12'h777;
rom[551] = 12'hccc;
rom[552] = 12'hccc;
rom[553] = 12'hccc;
rom[554] = 12'hccc;
rom[555] = 12'hccc;
rom[556] = 12'hccc;
rom[557] = 12'hccc;
rom[558] = 12'hccc;
rom[559] = 12'hccc;
rom[560] = 12'hccc;
rom[561] = 12'hccc;
rom[562] = 12'hccc;
rom[563] = 12'hccc;
rom[564] = 12'hccc;
rom[565] = 12'hccc;
rom[566] = 12'hccc;
rom[567] = 12'hccc;
rom[568] = 12'hccc;
rom[569] = 12'hccc;
rom[570] = 12'hccc;
rom[571] = 12'hccc;
rom[572] = 12'hccc;
rom[573] = 12'hccc;
rom[574] = 12'h777;
rom[575] = 12'h777;
rom[576] = 12'hccc;
rom[577] = 12'hccc;
rom[578] = 12'hccc;
rom[579] = 12'hccc;
rom[580] = 12'hccc;
rom[581] = 12'hccc;
rom[582] = 12'hccc;
rom[583] = 12'hccc;
rom[584] = 12'hccc;
rom[585] = 12'hccc;
rom[586] = 12'hccc;
rom[587] = 12'hccc;
rom[588] = 12'hccc;
rom[589] = 12'hccc;
rom[590] = 12'hccc;
rom[591] = 12'hccc;
rom[592] = 12'hccc;
rom[593] = 12'hccc;
rom[594] = 12'hccc;
rom[595] = 12'hccc;
rom[596] = 12'hccc;
rom[597] = 12'hccc;
rom[598] = 12'hccc;
rom[599] = 12'h777;
rom[600] = 12'h777;
rom[601] = 12'h777;
rom[602] = 12'h777;
rom[603] = 12'h777;
rom[604] = 12'h777;
rom[605] = 12'h777;
rom[606] = 12'h777;
rom[607] = 12'h777;
rom[608] = 12'h777;
rom[609] = 12'h777;
rom[610] = 12'h777;
rom[611] = 12'h777;
rom[612] = 12'h777;
rom[613] = 12'h777;
rom[614] = 12'h777;
rom[615] = 12'h777;
rom[616] = 12'h777;
rom[617] = 12'h777;
rom[618] = 12'h777;
rom[619] = 12'h777;
rom[620] = 12'h777;
rom[621] = 12'h777;
rom[622] = 12'h777;
rom[623] = 12'h777;
rom[624] = 12'h777;
  end
  endmodule

  module tile_eight_rom (                       //клетка с восьмёркой
  input  wire    [13:0]     addr,
  output wire    [11:0]     word
);

  logic [11:0] rom [(25 * 25)];

  assign word = rom[addr];

  initial begin
rom[0] = 12'h777;
rom[1] = 12'h777;
rom[2] = 12'h777;
rom[3] = 12'h777;
rom[4] = 12'h777;
rom[5] = 12'h777;
rom[6] = 12'h777;
rom[7] = 12'h777;
rom[8] = 12'h777;
rom[9] = 12'h777;
rom[10] = 12'h777;
rom[11] = 12'h777;
rom[12] = 12'h777;
rom[13] = 12'h777;
rom[14] = 12'h777;
rom[15] = 12'h777;
rom[16] = 12'h777;
rom[17] = 12'h777;
rom[18] = 12'h777;
rom[19] = 12'h777;
rom[20] = 12'h777;
rom[21] = 12'h777;
rom[22] = 12'h777;
rom[23] = 12'h777;
rom[24] = 12'h777;
rom[25] = 12'h777;
rom[26] = 12'hccc;
rom[27] = 12'hccc;
rom[28] = 12'hccc;
rom[29] = 12'hccc;
rom[30] = 12'hccc;
rom[31] = 12'hccc;
rom[32] = 12'hccc;
rom[33] = 12'hccc;
rom[34] = 12'hccc;
rom[35] = 12'hccc;
rom[36] = 12'hccc;
rom[37] = 12'hccc;
rom[38] = 12'hccc;
rom[39] = 12'hccc;
rom[40] = 12'hccc;
rom[41] = 12'hccc;
rom[42] = 12'hccc;
rom[43] = 12'hccc;
rom[44] = 12'hccc;
rom[45] = 12'hccc;
rom[46] = 12'hccc;
rom[47] = 12'hccc;
rom[48] = 12'hccc;
rom[49] = 12'h777;
rom[50] = 12'h777;
rom[51] = 12'hccc;
rom[52] = 12'hccc;
rom[53] = 12'hccc;
rom[54] = 12'hccc;
rom[55] = 12'hccc;
rom[56] = 12'hccc;
rom[57] = 12'hccc;
rom[58] = 12'hccc;
rom[59] = 12'hccc;
rom[60] = 12'hccc;
rom[61] = 12'hccc;
rom[62] = 12'hccc;
rom[63] = 12'hccc;
rom[64] = 12'hccc;
rom[65] = 12'hccc;
rom[66] = 12'hccc;
rom[67] = 12'hccc;
rom[68] = 12'hccc;
rom[69] = 12'hccc;
rom[70] = 12'hccc;
rom[71] = 12'hccc;
rom[72] = 12'hccc;
rom[73] = 12'hccc;
rom[74] = 12'h777;
rom[75] = 12'h777;
rom[76] = 12'hccc;
rom[77] = 12'hccc;
rom[78] = 12'hccc;
rom[79] = 12'hccc;
rom[80] = 12'hccc;
rom[81] = 12'hccc;
rom[82] = 12'hccc;
rom[83] = 12'hccc;
rom[84] = 12'hccc;
rom[85] = 12'hccc;
rom[86] = 12'hccc;
rom[87] = 12'hccc;
rom[88] = 12'hccc;
rom[89] = 12'hccc;
rom[90] = 12'hccc;
rom[91] = 12'hccc;
rom[92] = 12'hccc;
rom[93] = 12'hccc;
rom[94] = 12'hccc;
rom[95] = 12'hccc;
rom[96] = 12'hccc;
rom[97] = 12'hccc;
rom[98] = 12'hccc;
rom[99] = 12'h777;
rom[100] = 12'h777;
rom[101] = 12'hccc;
rom[102] = 12'hccc;
rom[103] = 12'hccc;
rom[104] = 12'hccc;
rom[105] = 12'hccc;
rom[106] = 12'hccc;
rom[107] = 12'hccc;
rom[108] = 12'hccc;
rom[109] = 12'hccc;
rom[110] = 12'hccc;
rom[111] = 12'hccc;
rom[112] = 12'hccc;
rom[113] = 12'hccc;
rom[114] = 12'hccc;
rom[115] = 12'hccc;
rom[116] = 12'hccc;
rom[117] = 12'hccc;
rom[118] = 12'hccc;
rom[119] = 12'hccc;
rom[120] = 12'hccc;
rom[121] = 12'hccc;
rom[122] = 12'hccc;
rom[123] = 12'hccc;
rom[124] = 12'h777;
rom[125] = 12'h777;
rom[126] = 12'hccc;
rom[127] = 12'hccc;
rom[128] = 12'hccc;
rom[129] = 12'hccc;
rom[130] = 12'hccc;
rom[131] = 12'hccc;
rom[132] = 12'hccc;
rom[133] = 12'hccc;
rom[134] = 12'hccc;
rom[135] = 12'hccc;
rom[136] = 12'hccc;
rom[137] = 12'hccc;
rom[138] = 12'hccc;
rom[139] = 12'hccc;
rom[140] = 12'hccc;
rom[141] = 12'hccc;
rom[142] = 12'hccc;
rom[143] = 12'hccc;
rom[144] = 12'hccc;
rom[145] = 12'hccc;
rom[146] = 12'hccc;
rom[147] = 12'hccc;
rom[148] = 12'hccc;
rom[149] = 12'h777;
rom[150] = 12'h777;
rom[151] = 12'hccc;
rom[152] = 12'hccc;
rom[153] = 12'hccc;
rom[154] = 12'hccc;
rom[155] = 12'hccc;
rom[156] = 12'hccc;
rom[157] = 12'hccc;
rom[158] = 12'hccc;
rom[159] = 12'hccc;
rom[160] = 12'hccc;
rom[161] = 12'hccc;
rom[162] = 12'hccc;
rom[163] = 12'hccc;
rom[164] = 12'hccc;
rom[165] = 12'hccc;
rom[166] = 12'hccc;
rom[167] = 12'hccc;
rom[168] = 12'hccc;
rom[169] = 12'hccc;
rom[170] = 12'hccc;
rom[171] = 12'hccc;
rom[172] = 12'hccc;
rom[173] = 12'hccc;
rom[174] = 12'h777;
rom[175] = 12'h777;
rom[176] = 12'hccc;
rom[177] = 12'hccc;
rom[178] = 12'hccc;
rom[179] = 12'hccc;
rom[180] = 12'hccc;
rom[181] = 12'hccc;
rom[182] = 12'hccc;
rom[183] = 12'hccc;
rom[184] = 12'h777;
rom[185] = 12'h777;
rom[186] = 12'h777;
rom[187] = 12'h777;
rom[188] = 12'h777;
rom[189] = 12'h777;
rom[190] = 12'h777;
rom[191] = 12'h777;
rom[192] = 12'hccc;
rom[193] = 12'hccc;
rom[194] = 12'hccc;
rom[195] = 12'hccc;
rom[196] = 12'hccc;
rom[197] = 12'hccc;
rom[198] = 12'hccc;
rom[199] = 12'h777;
rom[200] = 12'h777;
rom[201] = 12'hccc;
rom[202] = 12'hccc;
rom[203] = 12'hccc;
rom[204] = 12'hccc;
rom[205] = 12'hccc;
rom[206] = 12'hccc;
rom[207] = 12'hccc;
rom[208] = 12'h777;
rom[209] = 12'h777;
rom[210] = 12'h777;
rom[211] = 12'h777;
rom[212] = 12'h777;
rom[213] = 12'h777;
rom[214] = 12'h777;
rom[215] = 12'h777;
rom[216] = 12'h777;
rom[217] = 12'h777;
rom[218] = 12'hccc;
rom[219] = 12'hccc;
rom[220] = 12'hccc;
rom[221] = 12'hccc;
rom[222] = 12'hccc;
rom[223] = 12'hccc;
rom[224] = 12'h777;
rom[225] = 12'h777;
rom[226] = 12'hccc;
rom[227] = 12'hccc;
rom[228] = 12'hccc;
rom[229] = 12'hccc;
rom[230] = 12'hccc;
rom[231] = 12'hccc;
rom[232] = 12'hccc;
rom[233] = 12'h777;
rom[234] = 12'h777;
rom[235] = 12'h777;
rom[236] = 12'hccc;
rom[237] = 12'hccc;
rom[238] = 12'hccc;
rom[239] = 12'hccc;
rom[240] = 12'h777;
rom[241] = 12'h777;
rom[242] = 12'h777;
rom[243] = 12'hccc;
rom[244] = 12'hccc;
rom[245] = 12'hccc;
rom[246] = 12'hccc;
rom[247] = 12'hccc;
rom[248] = 12'hccc;
rom[249] = 12'h777;
rom[250] = 12'h777;
rom[251] = 12'hccc;
rom[252] = 12'hccc;
rom[253] = 12'hccc;
rom[254] = 12'hccc;
rom[255] = 12'hccc;
rom[256] = 12'hccc;
rom[257] = 12'hccc;
rom[258] = 12'h777;
rom[259] = 12'h777;
rom[260] = 12'h777;
rom[261] = 12'hccc;
rom[262] = 12'hccc;
rom[263] = 12'hccc;
rom[264] = 12'hccc;
rom[265] = 12'h777;
rom[266] = 12'h777;
rom[267] = 12'h777;
rom[268] = 12'hccc;
rom[269] = 12'hccc;
rom[270] = 12'hccc;
rom[271] = 12'hccc;
rom[272] = 12'hccc;
rom[273] = 12'hccc;
rom[274] = 12'h777;
rom[275] = 12'h777;
rom[276] = 12'hccc;
rom[277] = 12'hccc;
rom[278] = 12'hccc;
rom[279] = 12'hccc;
rom[280] = 12'hccc;
rom[281] = 12'hccc;
rom[282] = 12'hccc;
rom[283] = 12'hccc;
rom[284] = 12'h777;
rom[285] = 12'h777;
rom[286] = 12'h777;
rom[287] = 12'h777;
rom[288] = 12'h777;
rom[289] = 12'h777;
rom[290] = 12'h777;
rom[291] = 12'h777;
rom[292] = 12'hccc;
rom[293] = 12'hccc;
rom[294] = 12'hccc;
rom[295] = 12'hccc;
rom[296] = 12'hccc;
rom[297] = 12'hccc;
rom[298] = 12'hccc;
rom[299] = 12'h777;
rom[300] = 12'h777;
rom[301] = 12'hccc;
rom[302] = 12'hccc;
rom[303] = 12'hccc;
rom[304] = 12'hccc;
rom[305] = 12'hccc;
rom[306] = 12'hccc;
rom[307] = 12'hccc;
rom[308] = 12'hccc;
rom[309] = 12'h777;
rom[310] = 12'h777;
rom[311] = 12'h777;
rom[312] = 12'h777;
rom[313] = 12'h777;
rom[314] = 12'h777;
rom[315] = 12'h777;
rom[316] = 12'h777;
rom[317] = 12'hccc;
rom[318] = 12'hccc;
rom[319] = 12'hccc;
rom[320] = 12'hccc;
rom[321] = 12'hccc;
rom[322] = 12'hccc;
rom[323] = 12'hccc;
rom[324] = 12'h777;
rom[325] = 12'h777;
rom[326] = 12'hccc;
rom[327] = 12'hccc;
rom[328] = 12'hccc;
rom[329] = 12'hccc;
rom[330] = 12'hccc;
rom[331] = 12'hccc;
rom[332] = 12'hccc;
rom[333] = 12'h777;
rom[334] = 12'h777;
rom[335] = 12'h777;
rom[336] = 12'hccc;
rom[337] = 12'hccc;
rom[338] = 12'hccc;
rom[339] = 12'hccc;
rom[340] = 12'h777;
rom[341] = 12'h777;
rom[342] = 12'h777;
rom[343] = 12'hccc;
rom[344] = 12'hccc;
rom[345] = 12'hccc;
rom[346] = 12'hccc;
rom[347] = 12'hccc;
rom[348] = 12'hccc;
rom[349] = 12'h777;
rom[350] = 12'h777;
rom[351] = 12'hccc;
rom[352] = 12'hccc;
rom[353] = 12'hccc;
rom[354] = 12'hccc;
rom[355] = 12'hccc;
rom[356] = 12'hccc;
rom[357] = 12'hccc;
rom[358] = 12'h777;
rom[359] = 12'h777;
rom[360] = 12'h777;
rom[361] = 12'hccc;
rom[362] = 12'hccc;
rom[363] = 12'hccc;
rom[364] = 12'hccc;
rom[365] = 12'h777;
rom[366] = 12'h777;
rom[367] = 12'h777;
rom[368] = 12'hccc;
rom[369] = 12'hccc;
rom[370] = 12'hccc;
rom[371] = 12'hccc;
rom[372] = 12'hccc;
rom[373] = 12'hccc;
rom[374] = 12'h777;
rom[375] = 12'h777;
rom[376] = 12'hccc;
rom[377] = 12'hccc;
rom[378] = 12'hccc;
rom[379] = 12'hccc;
rom[380] = 12'hccc;
rom[381] = 12'hccc;
rom[382] = 12'hccc;
rom[383] = 12'h777;
rom[384] = 12'h777;
rom[385] = 12'h777;
rom[386] = 12'h777;
rom[387] = 12'h777;
rom[388] = 12'h777;
rom[389] = 12'h777;
rom[390] = 12'h777;
rom[391] = 12'h777;
rom[392] = 12'h777;
rom[393] = 12'hccc;
rom[394] = 12'hccc;
rom[395] = 12'hccc;
rom[396] = 12'hccc;
rom[397] = 12'hccc;
rom[398] = 12'hccc;
rom[399] = 12'h777;
rom[400] = 12'h777;
rom[401] = 12'hccc;
rom[402] = 12'hccc;
rom[403] = 12'hccc;
rom[404] = 12'hccc;
rom[405] = 12'hccc;
rom[406] = 12'hccc;
rom[407] = 12'hccc;
rom[408] = 12'hccc;
rom[409] = 12'h777;
rom[410] = 12'h777;
rom[411] = 12'h777;
rom[412] = 12'h777;
rom[413] = 12'h777;
rom[414] = 12'h777;
rom[415] = 12'h777;
rom[416] = 12'h777;
rom[417] = 12'hccc;
rom[418] = 12'hccc;
rom[419] = 12'hccc;
rom[420] = 12'hccc;
rom[421] = 12'hccc;
rom[422] = 12'hccc;
rom[423] = 12'hccc;
rom[424] = 12'h777;
rom[425] = 12'h777;
rom[426] = 12'hccc;
rom[427] = 12'hccc;
rom[428] = 12'hccc;
rom[429] = 12'hccc;
rom[430] = 12'hccc;
rom[431] = 12'hccc;
rom[432] = 12'hccc;
rom[433] = 12'hccc;
rom[434] = 12'hccc;
rom[435] = 12'hccc;
rom[436] = 12'hccc;
rom[437] = 12'hccc;
rom[438] = 12'hccc;
rom[439] = 12'hccc;
rom[440] = 12'hbbb;
rom[441] = 12'hccc;
rom[442] = 12'hccc;
rom[443] = 12'hccc;
rom[444] = 12'hccc;
rom[445] = 12'hccc;
rom[446] = 12'hccc;
rom[447] = 12'hccc;
rom[448] = 12'hccc;
rom[449] = 12'h777;
rom[450] = 12'h777;
rom[451] = 12'hccc;
rom[452] = 12'hccc;
rom[453] = 12'hccc;
rom[454] = 12'hccc;
rom[455] = 12'hccc;
rom[456] = 12'hccc;
rom[457] = 12'hccc;
rom[458] = 12'hccc;
rom[459] = 12'hccc;
rom[460] = 12'hccc;
rom[461] = 12'hccc;
rom[462] = 12'hccc;
rom[463] = 12'hccc;
rom[464] = 12'hccc;
rom[465] = 12'hbbb;
rom[466] = 12'hccc;
rom[467] = 12'hccc;
rom[468] = 12'hccc;
rom[469] = 12'hccc;
rom[470] = 12'hccc;
rom[471] = 12'hccc;
rom[472] = 12'hccc;
rom[473] = 12'hccc;
rom[474] = 12'h777;
rom[475] = 12'h777;
rom[476] = 12'hccc;
rom[477] = 12'hccc;
rom[478] = 12'hccc;
rom[479] = 12'hccc;
rom[480] = 12'hccc;
rom[481] = 12'hccc;
rom[482] = 12'hccc;
rom[483] = 12'hccc;
rom[484] = 12'hccc;
rom[485] = 12'hccc;
rom[486] = 12'hccc;
rom[487] = 12'hccc;
rom[488] = 12'hccc;
rom[489] = 12'hccc;
rom[490] = 12'hccc;
rom[491] = 12'hccc;
rom[492] = 12'hccc;
rom[493] = 12'hccc;
rom[494] = 12'hccc;
rom[495] = 12'hccc;
rom[496] = 12'hccc;
rom[497] = 12'hccc;
rom[498] = 12'hccc;
rom[499] = 12'h777;
rom[500] = 12'h777;
rom[501] = 12'hccc;
rom[502] = 12'hccc;
rom[503] = 12'hccc;
rom[504] = 12'hccc;
rom[505] = 12'hccc;
rom[506] = 12'hccc;
rom[507] = 12'hccc;
rom[508] = 12'hccc;
rom[509] = 12'hccc;
rom[510] = 12'hccc;
rom[511] = 12'hccc;
rom[512] = 12'hccc;
rom[513] = 12'hccc;
rom[514] = 12'hccc;
rom[515] = 12'hccc;
rom[516] = 12'hccc;
rom[517] = 12'hccc;
rom[518] = 12'hccc;
rom[519] = 12'hccc;
rom[520] = 12'hccc;
rom[521] = 12'hccc;
rom[522] = 12'hccc;
rom[523] = 12'hccc;
rom[524] = 12'h777;
rom[525] = 12'h777;
rom[526] = 12'hccc;
rom[527] = 12'hccc;
rom[528] = 12'hccc;
rom[529] = 12'hccc;
rom[530] = 12'hccc;
rom[531] = 12'hccc;
rom[532] = 12'hccc;
rom[533] = 12'hccc;
rom[534] = 12'hccc;
rom[535] = 12'hccc;
rom[536] = 12'hccc;
rom[537] = 12'hccc;
rom[538] = 12'hccc;
rom[539] = 12'hccc;
rom[540] = 12'hccc;
rom[541] = 12'hccc;
rom[542] = 12'hccc;
rom[543] = 12'hccc;
rom[544] = 12'hccc;
rom[545] = 12'hccc;
rom[546] = 12'hccc;
rom[547] = 12'hccc;
rom[548] = 12'hccc;
rom[549] = 12'h777;
rom[550] = 12'h777;
rom[551] = 12'hccc;
rom[552] = 12'hccc;
rom[553] = 12'hccc;
rom[554] = 12'hccc;
rom[555] = 12'hccc;
rom[556] = 12'hccc;
rom[557] = 12'hccc;
rom[558] = 12'hccc;
rom[559] = 12'hccc;
rom[560] = 12'hccc;
rom[561] = 12'hccc;
rom[562] = 12'hccc;
rom[563] = 12'hccc;
rom[564] = 12'hccc;
rom[565] = 12'hccc;
rom[566] = 12'hccc;
rom[567] = 12'hccc;
rom[568] = 12'hccc;
rom[569] = 12'hccc;
rom[570] = 12'hccc;
rom[571] = 12'hccc;
rom[572] = 12'hccc;
rom[573] = 12'hccc;
rom[574] = 12'h777;
rom[575] = 12'h777;
rom[576] = 12'hccc;
rom[577] = 12'hccc;
rom[578] = 12'hccc;
rom[579] = 12'hccc;
rom[580] = 12'hccc;
rom[581] = 12'hccc;
rom[582] = 12'hccc;
rom[583] = 12'hccc;
rom[584] = 12'hccc;
rom[585] = 12'hccc;
rom[586] = 12'hccc;
rom[587] = 12'hccc;
rom[588] = 12'hccc;
rom[589] = 12'hccc;
rom[590] = 12'hccc;
rom[591] = 12'hccc;
rom[592] = 12'hccc;
rom[593] = 12'hccc;
rom[594] = 12'hccc;
rom[595] = 12'hccc;
rom[596] = 12'hccc;
rom[597] = 12'hccc;
rom[598] = 12'hccc;
rom[599] = 12'h777;
rom[600] = 12'h777;
rom[601] = 12'h777;
rom[602] = 12'h777;
rom[603] = 12'h777;
rom[604] = 12'h777;
rom[605] = 12'h777;
rom[606] = 12'h777;
rom[607] = 12'h777;
rom[608] = 12'h777;
rom[609] = 12'h777;
rom[610] = 12'h777;
rom[611] = 12'h777;
rom[612] = 12'h777;
rom[613] = 12'h777;
rom[614] = 12'h777;
rom[615] = 12'h777;
rom[616] = 12'h777;
rom[617] = 12'h777;
rom[618] = 12'h777;
rom[619] = 12'h777;
rom[620] = 12'h777;
rom[621] = 12'h777;
rom[622] = 12'h777;
rom[623] = 12'h777;
rom[624] = 12'h777;
  end
  endmodule

module mine_rom (                       //клетка с миной
  input  wire    [13:0]     addr,
  output wire    [11:0]     word
);

  logic [11:0] rom [(25 * 25)];

  assign word = rom[addr];

  initial begin
rom[0] = 12'h777;
rom[1] = 12'h777;
rom[2] = 12'h777;
rom[3] = 12'h777;
rom[4] = 12'h777;
rom[5] = 12'h777;
rom[6] = 12'h777;
rom[7] = 12'h777;
rom[8] = 12'h777;
rom[9] = 12'h777;
rom[10] = 12'h777;
rom[11] = 12'h777;
rom[12] = 12'h777;
rom[13] = 12'h777;
rom[14] = 12'h777;
rom[15] = 12'h777;
rom[16] = 12'h777;
rom[17] = 12'h777;
rom[18] = 12'h777;
rom[19] = 12'h777;
rom[20] = 12'h777;
rom[21] = 12'h777;
rom[22] = 12'h777;
rom[23] = 12'h777;
rom[24] = 12'h777;
rom[25] = 12'h777;
rom[26] = 12'hccc;
rom[27] = 12'hccc;
rom[28] = 12'hccc;
rom[29] = 12'hccc;
rom[30] = 12'hccc;
rom[31] = 12'hccc;
rom[32] = 12'hccc;
rom[33] = 12'hccc;
rom[34] = 12'hccc;
rom[35] = 12'hccc;
rom[36] = 12'hccc;
rom[37] = 12'hccc;
rom[38] = 12'hccc;
rom[39] = 12'hccc;
rom[40] = 12'hccc;
rom[41] = 12'hccc;
rom[42] = 12'hccc;
rom[43] = 12'hccc;
rom[44] = 12'hccc;
rom[45] = 12'hccc;
rom[46] = 12'hccc;
rom[47] = 12'hccc;
rom[48] = 12'hccc;
rom[49] = 12'h777;
rom[50] = 12'h777;
rom[51] = 12'hccc;
rom[52] = 12'hccc;
rom[53] = 12'hccc;
rom[54] = 12'hccc;
rom[55] = 12'hccc;
rom[56] = 12'hccc;
rom[57] = 12'hccc;
rom[58] = 12'hccc;
rom[59] = 12'hccc;
rom[60] = 12'hccc;
rom[61] = 12'hccc;
rom[62] = 12'hccc;
rom[63] = 12'hccc;
rom[64] = 12'hccc;
rom[65] = 12'hccc;
rom[66] = 12'hccc;
rom[67] = 12'hccc;
rom[68] = 12'hccc;
rom[69] = 12'hccc;
rom[70] = 12'hccc;
rom[71] = 12'hccc;
rom[72] = 12'hccc;
rom[73] = 12'hccc;
rom[74] = 12'h777;
rom[75] = 12'h777;
rom[76] = 12'hccc;
rom[77] = 12'hccc;
rom[78] = 12'hccc;
rom[79] = 12'hccc;
rom[80] = 12'hccc;
rom[81] = 12'hccc;
rom[82] = 12'hccc;
rom[83] = 12'hccc;
rom[84] = 12'hccc;
rom[85] = 12'hccc;
rom[86] = 12'hccc;
rom[87] = 12'hccc;
rom[88] = 12'hccc;
rom[89] = 12'hccc;
rom[90] = 12'hccc;
rom[91] = 12'hccc;
rom[92] = 12'hccc;
rom[93] = 12'hccc;
rom[94] = 12'hccc;
rom[95] = 12'hccc;
rom[96] = 12'hccc;
rom[97] = 12'hccc;
rom[98] = 12'hccc;
rom[99] = 12'h777;
rom[100] = 12'h777;
rom[101] = 12'hccc;
rom[102] = 12'hccc;
rom[103] = 12'hccc;
rom[104] = 12'hccc;
rom[105] = 12'hccc;
rom[106] = 12'hccc;
rom[107] = 12'hccc;
rom[108] = 12'hccc;
rom[109] = 12'hccc;
rom[110] = 12'hccc;
rom[111] = 12'hccc;
rom[112] = 12'hccc;
rom[113] = 12'hccc;
rom[114] = 12'hccc;
rom[115] = 12'hccc;
rom[116] = 12'hccc;
rom[117] = 12'hccc;
rom[118] = 12'hccc;
rom[119] = 12'hccc;
rom[120] = 12'hccc;
rom[121] = 12'hccc;
rom[122] = 12'hccc;
rom[123] = 12'hccc;
rom[124] = 12'h777;
rom[125] = 12'h777;
rom[126] = 12'hccc;
rom[127] = 12'hccc;
rom[128] = 12'hccc;
rom[129] = 12'hccc;
rom[130] = 12'hccc;
rom[131] = 12'hccc;
rom[132] = 12'hccc;
rom[133] = 12'hccc;
rom[134] = 12'hccc;
rom[135] = 12'hccc;
rom[136] = 12'hccc;
rom[137] = 12'hccc;
rom[138] = 12'hccc;
rom[139] = 12'hccc;
rom[140] = 12'hccc;
rom[141] = 12'hccc;
rom[142] = 12'hccc;
rom[143] = 12'hccc;
rom[144] = 12'hccc;
rom[145] = 12'hccc;
rom[146] = 12'hccc;
rom[147] = 12'hccc;
rom[148] = 12'hccc;
rom[149] = 12'h777;
rom[150] = 12'h777;
rom[151] = 12'hccc;
rom[152] = 12'hccc;
rom[153] = 12'hccc;
rom[154] = 12'hccc;
rom[155] = 12'hccc;
rom[156] = 12'hccc;
rom[157] = 12'hccc;
rom[158] = 12'hccc;
rom[159] = 12'hccc;
rom[160] = 12'hccc;
rom[161] = 12'hccc;
rom[162] = 12'h000;
rom[163] = 12'hccc;
rom[164] = 12'hccc;
rom[165] = 12'hccc;
rom[166] = 12'hccc;
rom[167] = 12'hccc;
rom[168] = 12'hccc;
rom[169] = 12'hccc;
rom[170] = 12'hccc;
rom[171] = 12'hccc;
rom[172] = 12'hccc;
rom[173] = 12'hccc;
rom[174] = 12'h777;
rom[175] = 12'h777;
rom[176] = 12'hccc;
rom[177] = 12'hccc;
rom[178] = 12'hccc;
rom[179] = 12'hccc;
rom[180] = 12'hccc;
rom[181] = 12'hccc;
rom[182] = 12'hccc;
rom[183] = 12'hccc;
rom[184] = 12'hccc;
rom[185] = 12'hccc;
rom[186] = 12'hccc;
rom[187] = 12'h000;
rom[188] = 12'hccc;
rom[189] = 12'hccc;
rom[190] = 12'hccc;
rom[191] = 12'hccc;
rom[192] = 12'hccc;
rom[193] = 12'hccc;
rom[194] = 12'hccc;
rom[195] = 12'hccc;
rom[196] = 12'hccc;
rom[197] = 12'hccc;
rom[198] = 12'hccc;
rom[199] = 12'h777;
rom[200] = 12'h777;
rom[201] = 12'hccc;
rom[202] = 12'hccc;
rom[203] = 12'hccc;
rom[204] = 12'hccc;
rom[205] = 12'hccc;
rom[206] = 12'hccc;
rom[207] = 12'hccc;
rom[208] = 12'h000;
rom[209] = 12'hccc;
rom[210] = 12'h000;
rom[211] = 12'h000;
rom[212] = 12'h000;
rom[213] = 12'h000;
rom[214] = 12'h000;
rom[215] = 12'hccc;
rom[216] = 12'h000;
rom[217] = 12'hccc;
rom[218] = 12'hccc;
rom[219] = 12'hccc;
rom[220] = 12'hccc;
rom[221] = 12'hccc;
rom[222] = 12'hccc;
rom[223] = 12'hccc;
rom[224] = 12'h777;
rom[225] = 12'h777;
rom[226] = 12'hccc;
rom[227] = 12'hccc;
rom[228] = 12'hccc;
rom[229] = 12'hccc;
rom[230] = 12'hccc;
rom[231] = 12'hccc;
rom[232] = 12'hccc;
rom[233] = 12'hccc;
rom[234] = 12'h000;
rom[235] = 12'h000;
rom[236] = 12'h000;
rom[237] = 12'h000;
rom[238] = 12'h000;
rom[239] = 12'h000;
rom[240] = 12'h000;
rom[241] = 12'hccc;
rom[242] = 12'hccc;
rom[243] = 12'hccc;
rom[244] = 12'hccc;
rom[245] = 12'hccc;
rom[246] = 12'hccc;
rom[247] = 12'hccc;
rom[248] = 12'hccc;
rom[249] = 12'h777;
rom[250] = 12'h777;
rom[251] = 12'hccc;
rom[252] = 12'hccc;
rom[253] = 12'hccc;
rom[254] = 12'hccc;
rom[255] = 12'hccc;
rom[256] = 12'hccc;
rom[257] = 12'hccc;
rom[258] = 12'h000;
rom[259] = 12'h000;
rom[260] = 12'hfff;
rom[261] = 12'hfff;
rom[262] = 12'h000;
rom[263] = 12'h000;
rom[264] = 12'h000;
rom[265] = 12'h000;
rom[266] = 12'h000;
rom[267] = 12'hccc;
rom[268] = 12'hccc;
rom[269] = 12'hccc;
rom[270] = 12'hccc;
rom[271] = 12'hccc;
rom[272] = 12'hccc;
rom[273] = 12'hccc;
rom[274] = 12'h777;
rom[275] = 12'h777;
rom[276] = 12'hccc;
rom[277] = 12'hccc;
rom[278] = 12'hccc;
rom[279] = 12'hccc;
rom[280] = 12'hccc;
rom[281] = 12'hccc;
rom[282] = 12'hccc;
rom[283] = 12'h000;
rom[284] = 12'h000;
rom[285] = 12'hfff;
rom[286] = 12'hfff;
rom[287] = 12'h000;
rom[288] = 12'h000;
rom[289] = 12'h000;
rom[290] = 12'h000;
rom[291] = 12'h000;
rom[292] = 12'hccc;
rom[293] = 12'hccc;
rom[294] = 12'hccc;
rom[295] = 12'hccc;
rom[296] = 12'hccc;
rom[297] = 12'hccc;
rom[298] = 12'hccc;
rom[299] = 12'h777;
rom[300] = 12'h777;
rom[301] = 12'hccc;
rom[302] = 12'hccc;
rom[303] = 12'hccc;
rom[304] = 12'hccc;
rom[305] = 12'hccc;
rom[306] = 12'h000;
rom[307] = 12'h000;
rom[308] = 12'h000;
rom[309] = 12'h000;
rom[310] = 12'h000;
rom[311] = 12'h000;
rom[312] = 12'h000;
rom[313] = 12'h000;
rom[314] = 12'h000;
rom[315] = 12'h000;
rom[316] = 12'h000;
rom[317] = 12'h000;
rom[318] = 12'h000;
rom[319] = 12'hccc;
rom[320] = 12'hccc;
rom[321] = 12'hccc;
rom[322] = 12'hccc;
rom[323] = 12'hccc;
rom[324] = 12'h777;
rom[325] = 12'h777;
rom[326] = 12'hccc;
rom[327] = 12'hccc;
rom[328] = 12'hccc;
rom[329] = 12'hccc;
rom[330] = 12'hccc;
rom[331] = 12'hccc;
rom[332] = 12'hccc;
rom[333] = 12'h000;
rom[334] = 12'h000;
rom[335] = 12'h000;
rom[336] = 12'h000;
rom[337] = 12'h000;
rom[338] = 12'h000;
rom[339] = 12'h000;
rom[340] = 12'h000;
rom[341] = 12'h000;
rom[342] = 12'hccc;
rom[343] = 12'hccc;
rom[344] = 12'hccc;
rom[345] = 12'hccc;
rom[346] = 12'hccc;
rom[347] = 12'hccc;
rom[348] = 12'hccc;
rom[349] = 12'h777;
rom[350] = 12'h777;
rom[351] = 12'hccc;
rom[352] = 12'hccc;
rom[353] = 12'hccc;
rom[354] = 12'hccc;
rom[355] = 12'hccc;
rom[356] = 12'hccc;
rom[357] = 12'hccc;
rom[358] = 12'h000;
rom[359] = 12'h000;
rom[360] = 12'h000;
rom[361] = 12'h000;
rom[362] = 12'h000;
rom[363] = 12'h000;
rom[364] = 12'h000;
rom[365] = 12'h000;
rom[366] = 12'h000;
rom[367] = 12'hccc;
rom[368] = 12'hccc;
rom[369] = 12'hccc;
rom[370] = 12'hccc;
rom[371] = 12'hccc;
rom[372] = 12'hccc;
rom[373] = 12'hccc;
rom[374] = 12'h777;
rom[375] = 12'h777;
rom[376] = 12'hccc;
rom[377] = 12'hccc;
rom[378] = 12'hccc;
rom[379] = 12'hccc;
rom[380] = 12'hccc;
rom[381] = 12'hccc;
rom[382] = 12'hccc;
rom[383] = 12'hccc;
rom[384] = 12'h000;
rom[385] = 12'h000;
rom[386] = 12'h000;
rom[387] = 12'h000;
rom[388] = 12'h000;
rom[389] = 12'h000;
rom[390] = 12'h000;
rom[391] = 12'hccc;
rom[392] = 12'hccc;
rom[393] = 12'hccc;
rom[394] = 12'hccc;
rom[395] = 12'hccc;
rom[396] = 12'hccc;
rom[397] = 12'hccc;
rom[398] = 12'hccc;
rom[399] = 12'h777;
rom[400] = 12'h777;
rom[401] = 12'hccc;
rom[402] = 12'hccc;
rom[403] = 12'hccc;
rom[404] = 12'hccc;
rom[405] = 12'hccc;
rom[406] = 12'hccc;
rom[407] = 12'hccc;
rom[408] = 12'h000;
rom[409] = 12'hccc;
rom[410] = 12'h000;
rom[411] = 12'h000;
rom[412] = 12'h000;
rom[413] = 12'h000;
rom[414] = 12'h000;
rom[415] = 12'hccc;
rom[416] = 12'h000;
rom[417] = 12'hccc;
rom[418] = 12'hccc;
rom[419] = 12'hccc;
rom[420] = 12'hccc;
rom[421] = 12'hccc;
rom[422] = 12'hccc;
rom[423] = 12'hccc;
rom[424] = 12'h777;
rom[425] = 12'h777;
rom[426] = 12'hccc;
rom[427] = 12'hccc;
rom[428] = 12'hccc;
rom[429] = 12'hccc;
rom[430] = 12'hccc;
rom[431] = 12'hccc;
rom[432] = 12'hccc;
rom[433] = 12'hccc;
rom[434] = 12'hccc;
rom[435] = 12'hccc;
rom[436] = 12'hccc;
rom[437] = 12'h000;
rom[438] = 12'hccc;
rom[439] = 12'hccc;
rom[440] = 12'hbbb;
rom[441] = 12'hccc;
rom[442] = 12'hccc;
rom[443] = 12'hccc;
rom[444] = 12'hccc;
rom[445] = 12'hccc;
rom[446] = 12'hccc;
rom[447] = 12'hccc;
rom[448] = 12'hccc;
rom[449] = 12'h777;
rom[450] = 12'h777;
rom[451] = 12'hccc;
rom[452] = 12'hccc;
rom[453] = 12'hccc;
rom[454] = 12'hccc;
rom[455] = 12'hccc;
rom[456] = 12'hccc;
rom[457] = 12'hccc;
rom[458] = 12'hccc;
rom[459] = 12'hccc;
rom[460] = 12'hccc;
rom[461] = 12'hccc;
rom[462] = 12'h000;
rom[463] = 12'hccc;
rom[464] = 12'hccc;
rom[465] = 12'hbbb;
rom[466] = 12'hccc;
rom[467] = 12'hccc;
rom[468] = 12'hccc;
rom[469] = 12'hccc;
rom[470] = 12'hccc;
rom[471] = 12'hccc;
rom[472] = 12'hccc;
rom[473] = 12'hccc;
rom[474] = 12'h777;
rom[475] = 12'h777;
rom[476] = 12'hccc;
rom[477] = 12'hccc;
rom[478] = 12'hccc;
rom[479] = 12'hccc;
rom[480] = 12'hccc;
rom[481] = 12'hccc;
rom[482] = 12'hccc;
rom[483] = 12'hccc;
rom[484] = 12'hccc;
rom[485] = 12'hccc;
rom[486] = 12'hccc;
rom[487] = 12'hccc;
rom[488] = 12'hccc;
rom[489] = 12'hccc;
rom[490] = 12'hccc;
rom[491] = 12'hccc;
rom[492] = 12'hccc;
rom[493] = 12'hccc;
rom[494] = 12'hccc;
rom[495] = 12'hccc;
rom[496] = 12'hccc;
rom[497] = 12'hccc;
rom[498] = 12'hccc;
rom[499] = 12'h777;
rom[500] = 12'h777;
rom[501] = 12'hccc;
rom[502] = 12'hccc;
rom[503] = 12'hccc;
rom[504] = 12'hccc;
rom[505] = 12'hccc;
rom[506] = 12'hccc;
rom[507] = 12'hccc;
rom[508] = 12'hccc;
rom[509] = 12'hccc;
rom[510] = 12'hccc;
rom[511] = 12'hccc;
rom[512] = 12'hccc;
rom[513] = 12'hccc;
rom[514] = 12'hccc;
rom[515] = 12'hccc;
rom[516] = 12'hccc;
rom[517] = 12'hccc;
rom[518] = 12'hccc;
rom[519] = 12'hccc;
rom[520] = 12'hccc;
rom[521] = 12'hccc;
rom[522] = 12'hccc;
rom[523] = 12'hccc;
rom[524] = 12'h777;
rom[525] = 12'h777;
rom[526] = 12'hccc;
rom[527] = 12'hccc;
rom[528] = 12'hccc;
rom[529] = 12'hccc;
rom[530] = 12'hccc;
rom[531] = 12'hccc;
rom[532] = 12'hccc;
rom[533] = 12'hccc;
rom[534] = 12'hccc;
rom[535] = 12'hccc;
rom[536] = 12'hccc;
rom[537] = 12'hccc;
rom[538] = 12'hccc;
rom[539] = 12'hccc;
rom[540] = 12'hccc;
rom[541] = 12'hccc;
rom[542] = 12'hccc;
rom[543] = 12'hccc;
rom[544] = 12'hccc;
rom[545] = 12'hccc;
rom[546] = 12'hccc;
rom[547] = 12'hccc;
rom[548] = 12'hccc;
rom[549] = 12'h777;
rom[550] = 12'h777;
rom[551] = 12'hccc;
rom[552] = 12'hccc;
rom[553] = 12'hccc;
rom[554] = 12'hccc;
rom[555] = 12'hccc;
rom[556] = 12'hccc;
rom[557] = 12'hccc;
rom[558] = 12'hccc;
rom[559] = 12'hccc;
rom[560] = 12'hccc;
rom[561] = 12'hccc;
rom[562] = 12'hccc;
rom[563] = 12'hccc;
rom[564] = 12'hccc;
rom[565] = 12'hccc;
rom[566] = 12'hccc;
rom[567] = 12'hccc;
rom[568] = 12'hccc;
rom[569] = 12'hccc;
rom[570] = 12'hccc;
rom[571] = 12'hccc;
rom[572] = 12'hccc;
rom[573] = 12'hccc;
rom[574] = 12'h777;
rom[575] = 12'h777;
rom[576] = 12'hccc;
rom[577] = 12'hccc;
rom[578] = 12'hccc;
rom[579] = 12'hccc;
rom[580] = 12'hccc;
rom[581] = 12'hccc;
rom[582] = 12'hccc;
rom[583] = 12'hccc;
rom[584] = 12'hccc;
rom[585] = 12'hccc;
rom[586] = 12'hccc;
rom[587] = 12'hccc;
rom[588] = 12'hccc;
rom[589] = 12'hccc;
rom[590] = 12'hccc;
rom[591] = 12'hccc;
rom[592] = 12'hccc;
rom[593] = 12'hccc;
rom[594] = 12'hccc;
rom[595] = 12'hccc;
rom[596] = 12'hccc;
rom[597] = 12'hccc;
rom[598] = 12'hccc;
rom[599] = 12'h777;
rom[600] = 12'h777;
rom[601] = 12'h777;
rom[602] = 12'h777;
rom[603] = 12'h777;
rom[604] = 12'h777;
rom[605] = 12'h777;
rom[606] = 12'h777;
rom[607] = 12'h777;
rom[608] = 12'h777;
rom[609] = 12'h777;
rom[610] = 12'h777;
rom[611] = 12'h777;
rom[612] = 12'h777;
rom[613] = 12'h777;
rom[614] = 12'h777;
rom[615] = 12'h777;
rom[616] = 12'h777;
rom[617] = 12'h777;
rom[618] = 12'h777;
rom[619] = 12'h777;
rom[620] = 12'h777;
rom[621] = 12'h777;
rom[622] = 12'h777;
rom[623] = 12'h777;
rom[624] = 12'h777;
  end
  endmodule

module mine_exp_rom (                       //клетка с миной взрыв
  input  wire    [13:0]     addr,
  output wire    [11:0]     word
);

  logic [11:0] rom [(25 * 25)];

  assign word = rom[addr];

  initial begin
rom[0] = 12'h777;
rom[1] = 12'h777;
rom[2] = 12'h777;
rom[3] = 12'h777;
rom[4] = 12'h777;
rom[5] = 12'h777;
rom[6] = 12'h777;
rom[7] = 12'h777;
rom[8] = 12'h777;
rom[9] = 12'h777;
rom[10] = 12'h777;
rom[11] = 12'h777;
rom[12] = 12'h777;
rom[13] = 12'h777;
rom[14] = 12'h777;
rom[15] = 12'h777;
rom[16] = 12'h777;
rom[17] = 12'h777;
rom[18] = 12'h777;
rom[19] = 12'h777;
rom[20] = 12'h777;
rom[21] = 12'h777;
rom[22] = 12'h777;
rom[23] = 12'h777;
rom[24] = 12'h777;
rom[25] = 12'h777;
rom[26] = 12'h00f;
rom[27] = 12'h00f;
rom[28] = 12'h00f;
rom[29] = 12'h00f;
rom[30] = 12'h00f;
rom[31] = 12'h00f;
rom[32] = 12'h00f;
rom[33] = 12'h00f;
rom[34] = 12'h00f;
rom[35] = 12'h00f;
rom[36] = 12'h00f;
rom[37] = 12'h00f;
rom[38] = 12'h00f;
rom[39] = 12'h00f;
rom[40] = 12'h00f;
rom[41] = 12'h00f;
rom[42] = 12'h00f;
rom[43] = 12'h00f;
rom[44] = 12'h00f;
rom[45] = 12'h00f;
rom[46] = 12'h00f;
rom[47] = 12'h00f;
rom[48] = 12'h00f;
rom[49] = 12'h777;
rom[50] = 12'h777;
rom[51] = 12'h00f;
rom[52] = 12'h00f;
rom[53] = 12'h00f;
rom[54] = 12'h00f;
rom[55] = 12'h00f;
rom[56] = 12'h00f;
rom[57] = 12'h00f;
rom[58] = 12'h00f;
rom[59] = 12'h00f;
rom[60] = 12'h00f;
rom[61] = 12'h00f;
rom[62] = 12'h00f;
rom[63] = 12'h00f;
rom[64] = 12'h00f;
rom[65] = 12'h00f;
rom[66] = 12'h00f;
rom[67] = 12'h00f;
rom[68] = 12'h00f;
rom[69] = 12'h00f;
rom[70] = 12'h00f;
rom[71] = 12'h00f;
rom[72] = 12'h00f;
rom[73] = 12'h00f;
rom[74] = 12'h777;
rom[75] = 12'h777;
rom[76] = 12'h00f;
rom[77] = 12'h00f;
rom[78] = 12'h00f;
rom[79] = 12'h00f;
rom[80] = 12'h00f;
rom[81] = 12'h00f;
rom[82] = 12'h00f;
rom[83] = 12'h00f;
rom[84] = 12'h00f;
rom[85] = 12'h00f;
rom[86] = 12'h00f;
rom[87] = 12'h00f;
rom[88] = 12'h00f;
rom[89] = 12'h00f;
rom[90] = 12'h00f;
rom[91] = 12'h00f;
rom[92] = 12'h00f;
rom[93] = 12'h00f;
rom[94] = 12'h00f;
rom[95] = 12'h00f;
rom[96] = 12'h00f;
rom[97] = 12'h00f;
rom[98] = 12'h00f;
rom[99] = 12'h777;
rom[100] = 12'h777;
rom[101] = 12'h00f;
rom[102] = 12'h00f;
rom[103] = 12'h00f;
rom[104] = 12'h00f;
rom[105] = 12'h00f;
rom[106] = 12'h00f;
rom[107] = 12'h00f;
rom[108] = 12'h00f;
rom[109] = 12'h00f;
rom[110] = 12'h00f;
rom[111] = 12'h00f;
rom[112] = 12'h00f;
rom[113] = 12'h00f;
rom[114] = 12'h00f;
rom[115] = 12'h00f;
rom[116] = 12'h00f;
rom[117] = 12'h00f;
rom[118] = 12'h00f;
rom[119] = 12'h00f;
rom[120] = 12'h00f;
rom[121] = 12'h00f;
rom[122] = 12'h00f;
rom[123] = 12'h00f;
rom[124] = 12'h777;
rom[125] = 12'h777;
rom[126] = 12'h00f;
rom[127] = 12'h00f;
rom[128] = 12'h00f;
rom[129] = 12'h00f;
rom[130] = 12'h00f;
rom[131] = 12'h00f;
rom[132] = 12'h00f;
rom[133] = 12'h00f;
rom[134] = 12'h00f;
rom[135] = 12'h00f;
rom[136] = 12'h00f;
rom[137] = 12'h00f;
rom[138] = 12'h00f;
rom[139] = 12'h00f;
rom[140] = 12'h00f;
rom[141] = 12'h00f;
rom[142] = 12'h00f;
rom[143] = 12'h00f;
rom[144] = 12'h00f;
rom[145] = 12'h00f;
rom[146] = 12'h00f;
rom[147] = 12'h00f;
rom[148] = 12'h00f;
rom[149] = 12'h777;
rom[150] = 12'h777;
rom[151] = 12'h00f;
rom[152] = 12'h00f;
rom[153] = 12'h00f;
rom[154] = 12'h00f;
rom[155] = 12'h00f;
rom[156] = 12'h00f;
rom[157] = 12'h00f;
rom[158] = 12'h00f;
rom[159] = 12'h00f;
rom[160] = 12'h00f;
rom[161] = 12'h00f;
rom[162] = 12'h000;
rom[163] = 12'h00f;
rom[164] = 12'h00f;
rom[165] = 12'h00f;
rom[166] = 12'h00f;
rom[167] = 12'h00f;
rom[168] = 12'h00f;
rom[169] = 12'h00f;
rom[170] = 12'h00f;
rom[171] = 12'h00f;
rom[172] = 12'h00f;
rom[173] = 12'h00f;
rom[174] = 12'h777;
rom[175] = 12'h777;
rom[176] = 12'h00f;
rom[177] = 12'h00f;
rom[178] = 12'h00f;
rom[179] = 12'h00f;
rom[180] = 12'h00f;
rom[181] = 12'h00f;
rom[182] = 12'h00f;
rom[183] = 12'h00f;
rom[184] = 12'h00f;
rom[185] = 12'h00f;
rom[186] = 12'h00f;
rom[187] = 12'h000;
rom[188] = 12'h00f;
rom[189] = 12'h00f;
rom[190] = 12'h00f;
rom[191] = 12'h00f;
rom[192] = 12'h00f;
rom[193] = 12'h00f;
rom[194] = 12'h00f;
rom[195] = 12'h00f;
rom[196] = 12'h00f;
rom[197] = 12'h00f;
rom[198] = 12'h00f;
rom[199] = 12'h777;
rom[200] = 12'h777;
rom[201] = 12'h00f;
rom[202] = 12'h00f;
rom[203] = 12'h00f;
rom[204] = 12'h00f;
rom[205] = 12'h00f;
rom[206] = 12'h00f;
rom[207] = 12'h00f;
rom[208] = 12'h000;
rom[209] = 12'h00f;
rom[210] = 12'h000;
rom[211] = 12'h000;
rom[212] = 12'h000;
rom[213] = 12'h000;
rom[214] = 12'h000;
rom[215] = 12'h00f;
rom[216] = 12'h000;
rom[217] = 12'h00f;
rom[218] = 12'h00f;
rom[219] = 12'h00f;
rom[220] = 12'h00f;
rom[221] = 12'h00f;
rom[222] = 12'h00f;
rom[223] = 12'h00f;
rom[224] = 12'h777;
rom[225] = 12'h777;
rom[226] = 12'h00f;
rom[227] = 12'h00f;
rom[228] = 12'h00f;
rom[229] = 12'h00f;
rom[230] = 12'h00f;
rom[231] = 12'h00f;
rom[232] = 12'h00f;
rom[233] = 12'h00f;
rom[234] = 12'h000;
rom[235] = 12'h000;
rom[236] = 12'h000;
rom[237] = 12'h000;
rom[238] = 12'h000;
rom[239] = 12'h000;
rom[240] = 12'h000;
rom[241] = 12'h00f;
rom[242] = 12'h00f;
rom[243] = 12'h00f;
rom[244] = 12'h00f;
rom[245] = 12'h00f;
rom[246] = 12'h00f;
rom[247] = 12'h00f;
rom[248] = 12'h00f;
rom[249] = 12'h777;
rom[250] = 12'h777;
rom[251] = 12'h00f;
rom[252] = 12'h00f;
rom[253] = 12'h00f;
rom[254] = 12'h00f;
rom[255] = 12'h00f;
rom[256] = 12'h00f;
rom[257] = 12'h00f;
rom[258] = 12'h000;
rom[259] = 12'h000;
rom[260] = 12'hfff;
rom[261] = 12'hfff;
rom[262] = 12'h000;
rom[263] = 12'h000;
rom[264] = 12'h000;
rom[265] = 12'h000;
rom[266] = 12'h000;
rom[267] = 12'h00f;
rom[268] = 12'h00f;
rom[269] = 12'h00f;
rom[270] = 12'h00f;
rom[271] = 12'h00f;
rom[272] = 12'h00f;
rom[273] = 12'h00f;
rom[274] = 12'h777;
rom[275] = 12'h777;
rom[276] = 12'h00f;
rom[277] = 12'h00f;
rom[278] = 12'h00f;
rom[279] = 12'h00f;
rom[280] = 12'h00f;
rom[281] = 12'h00f;
rom[282] = 12'h00f;
rom[283] = 12'h000;
rom[284] = 12'h000;
rom[285] = 12'hfff;
rom[286] = 12'hfff;
rom[287] = 12'h000;
rom[288] = 12'h000;
rom[289] = 12'h000;
rom[290] = 12'h000;
rom[291] = 12'h000;
rom[292] = 12'h00f;
rom[293] = 12'h00f;
rom[294] = 12'h00f;
rom[295] = 12'h00f;
rom[296] = 12'h00f;
rom[297] = 12'h00f;
rom[298] = 12'h00f;
rom[299] = 12'h777;
rom[300] = 12'h777;
rom[301] = 12'h00f;
rom[302] = 12'h00f;
rom[303] = 12'h00f;
rom[304] = 12'h00f;
rom[305] = 12'h00f;
rom[306] = 12'h000;
rom[307] = 12'h000;
rom[308] = 12'h000;
rom[309] = 12'h000;
rom[310] = 12'h000;
rom[311] = 12'h000;
rom[312] = 12'h000;
rom[313] = 12'h000;
rom[314] = 12'h000;
rom[315] = 12'h000;
rom[316] = 12'h000;
rom[317] = 12'h000;
rom[318] = 12'h000;
rom[319] = 12'h00f;
rom[320] = 12'h00f;
rom[321] = 12'h00f;
rom[322] = 12'h00f;
rom[323] = 12'h00f;
rom[324] = 12'h777;
rom[325] = 12'h777;
rom[326] = 12'h00f;
rom[327] = 12'h00f;
rom[328] = 12'h00f;
rom[329] = 12'h00f;
rom[330] = 12'h00f;
rom[331] = 12'h00f;
rom[332] = 12'h00f;
rom[333] = 12'h000;
rom[334] = 12'h000;
rom[335] = 12'h000;
rom[336] = 12'h000;
rom[337] = 12'h000;
rom[338] = 12'h000;
rom[339] = 12'h000;
rom[340] = 12'h000;
rom[341] = 12'h000;
rom[342] = 12'h00f;
rom[343] = 12'h00f;
rom[344] = 12'h00f;
rom[345] = 12'h00f;
rom[346] = 12'h00f;
rom[347] = 12'h00f;
rom[348] = 12'h00f;
rom[349] = 12'h777;
rom[350] = 12'h777;
rom[351] = 12'h00f;
rom[352] = 12'h00f;
rom[353] = 12'h00f;
rom[354] = 12'h00f;
rom[355] = 12'h00f;
rom[356] = 12'h00f;
rom[357] = 12'h00f;
rom[358] = 12'h000;
rom[359] = 12'h000;
rom[360] = 12'h000;
rom[361] = 12'h000;
rom[362] = 12'h000;
rom[363] = 12'h000;
rom[364] = 12'h000;
rom[365] = 12'h000;
rom[366] = 12'h000;
rom[367] = 12'h00f;
rom[368] = 12'h00f;
rom[369] = 12'h00f;
rom[370] = 12'h00f;
rom[371] = 12'h00f;
rom[372] = 12'h00f;
rom[373] = 12'h00f;
rom[374] = 12'h777;
rom[375] = 12'h777;
rom[376] = 12'h00f;
rom[377] = 12'h00f;
rom[378] = 12'h00f;
rom[379] = 12'h00f;
rom[380] = 12'h00f;
rom[381] = 12'h00f;
rom[382] = 12'h00f;
rom[383] = 12'h00f;
rom[384] = 12'h000;
rom[385] = 12'h000;
rom[386] = 12'h000;
rom[387] = 12'h000;
rom[388] = 12'h000;
rom[389] = 12'h000;
rom[390] = 12'h000;
rom[391] = 12'h00f;
rom[392] = 12'h00f;
rom[393] = 12'h00f;
rom[394] = 12'h00f;
rom[395] = 12'h00f;
rom[396] = 12'h00f;
rom[397] = 12'h00f;
rom[398] = 12'h00f;
rom[399] = 12'h777;
rom[400] = 12'h777;
rom[401] = 12'h00f;
rom[402] = 12'h00f;
rom[403] = 12'h00f;
rom[404] = 12'h00f;
rom[405] = 12'h00f;
rom[406] = 12'h00f;
rom[407] = 12'h00f;
rom[408] = 12'h000;
rom[409] = 12'h00f;
rom[410] = 12'h000;
rom[411] = 12'h000;
rom[412] = 12'h000;
rom[413] = 12'h000;
rom[414] = 12'h000;
rom[415] = 12'h00f;
rom[416] = 12'h000;
rom[417] = 12'h00f;
rom[418] = 12'h00f;
rom[419] = 12'h00f;
rom[420] = 12'h00f;
rom[421] = 12'h00f;
rom[422] = 12'h00f;
rom[423] = 12'h00f;
rom[424] = 12'h777;
rom[425] = 12'h777;
rom[426] = 12'h00f;
rom[427] = 12'h00f;
rom[428] = 12'h00f;
rom[429] = 12'h00f;
rom[430] = 12'h00f;
rom[431] = 12'h00f;
rom[432] = 12'h00f;
rom[433] = 12'h00f;
rom[434] = 12'h00f;
rom[435] = 12'h00f;
rom[436] = 12'h00f;
rom[437] = 12'h000;
rom[438] = 12'h00f;
rom[439] = 12'h00f;
rom[440] = 12'h00f;
rom[441] = 12'h00f;
rom[442] = 12'h00f;
rom[443] = 12'h00f;
rom[444] = 12'h00f;
rom[445] = 12'h00f;
rom[446] = 12'h00f;
rom[447] = 12'h00f;
rom[448] = 12'h00f;
rom[449] = 12'h777;
rom[450] = 12'h777;
rom[451] = 12'h00f;
rom[452] = 12'h00f;
rom[453] = 12'h00f;
rom[454] = 12'h00f;
rom[455] = 12'h00f;
rom[456] = 12'h00f;
rom[457] = 12'h00f;
rom[458] = 12'h00f;
rom[459] = 12'h00f;
rom[460] = 12'h00f;
rom[461] = 12'h00f;
rom[462] = 12'h000;
rom[463] = 12'h00f;
rom[464] = 12'h00f;
rom[465] = 12'h00f;
rom[466] = 12'h00f;
rom[467] = 12'h00f;
rom[468] = 12'h00f;
rom[469] = 12'h00f;
rom[470] = 12'h00f;
rom[471] = 12'h00f;
rom[472] = 12'h00f;
rom[473] = 12'h00f;
rom[474] = 12'h777;
rom[475] = 12'h777;
rom[476] = 12'h00f;
rom[477] = 12'h00f;
rom[478] = 12'h00f;
rom[479] = 12'h00f;
rom[480] = 12'h00f;
rom[481] = 12'h00f;
rom[482] = 12'h00f;
rom[483] = 12'h00f;
rom[484] = 12'h00f;
rom[485] = 12'h00f;
rom[486] = 12'h00f;
rom[487] = 12'h00f;
rom[488] = 12'h00f;
rom[489] = 12'h00f;
rom[490] = 12'h00f;
rom[491] = 12'h00f;
rom[492] = 12'h00f;
rom[493] = 12'h00f;
rom[494] = 12'h00f;
rom[495] = 12'h00f;
rom[496] = 12'h00f;
rom[497] = 12'h00f;
rom[498] = 12'h00f;
rom[499] = 12'h777;
rom[500] = 12'h777;
rom[501] = 12'h00f;
rom[502] = 12'h00f;
rom[503] = 12'h00f;
rom[504] = 12'h00f;
rom[505] = 12'h00f;
rom[506] = 12'h00f;
rom[507] = 12'h00f;
rom[508] = 12'h00f;
rom[509] = 12'h00f;
rom[510] = 12'h00f;
rom[511] = 12'h00f;
rom[512] = 12'h00f;
rom[513] = 12'h00f;
rom[514] = 12'h00f;
rom[515] = 12'h00f;
rom[516] = 12'h00f;
rom[517] = 12'h00f;
rom[518] = 12'h00f;
rom[519] = 12'h00f;
rom[520] = 12'h00f;
rom[521] = 12'h00f;
rom[522] = 12'h00f;
rom[523] = 12'h00f;
rom[524] = 12'h777;
rom[525] = 12'h777;
rom[526] = 12'h00f;
rom[527] = 12'h00f;
rom[528] = 12'h00f;
rom[529] = 12'h00f;
rom[530] = 12'h00f;
rom[531] = 12'h00f;
rom[532] = 12'h00f;
rom[533] = 12'h00f;
rom[534] = 12'h00f;
rom[535] = 12'h00f;
rom[536] = 12'h00f;
rom[537] = 12'h00f;
rom[538] = 12'h00f;
rom[539] = 12'h00f;
rom[540] = 12'h00f;
rom[541] = 12'h00f;
rom[542] = 12'h00f;
rom[543] = 12'h00f;
rom[544] = 12'h00f;
rom[545] = 12'h00f;
rom[546] = 12'h00f;
rom[547] = 12'h00f;
rom[548] = 12'h00f;
rom[549] = 12'h777;
rom[550] = 12'h777;
rom[551] = 12'h00f;
rom[552] = 12'h00f;
rom[553] = 12'h00f;
rom[554] = 12'h00f;
rom[555] = 12'h00f;
rom[556] = 12'h00f;
rom[557] = 12'h00f;
rom[558] = 12'h00f;
rom[559] = 12'h00f;
rom[560] = 12'h00f;
rom[561] = 12'h00f;
rom[562] = 12'h00f;
rom[563] = 12'h00f;
rom[564] = 12'h00f;
rom[565] = 12'h00f;
rom[566] = 12'h00f;
rom[567] = 12'h00f;
rom[568] = 12'h00f;
rom[569] = 12'h00f;
rom[570] = 12'h00f;
rom[571] = 12'h00f;
rom[572] = 12'h00f;
rom[573] = 12'h00f;
rom[574] = 12'h777;
rom[575] = 12'h777;
rom[576] = 12'h00f;
rom[577] = 12'h00f;
rom[578] = 12'h00f;
rom[579] = 12'h00f;
rom[580] = 12'h00f;
rom[581] = 12'h00f;
rom[582] = 12'h00f;
rom[583] = 12'h00f;
rom[584] = 12'h00f;
rom[585] = 12'h00f;
rom[586] = 12'h00f;
rom[587] = 12'h00f;
rom[588] = 12'h00f;
rom[589] = 12'h00f;
rom[590] = 12'h00f;
rom[591] = 12'h00f;
rom[592] = 12'h00f;
rom[593] = 12'h00f;
rom[594] = 12'h00f;
rom[595] = 12'h00f;
rom[596] = 12'h00f;
rom[597] = 12'h00f;
rom[598] = 12'h00f;
rom[599] = 12'h777;
rom[600] = 12'h777;
rom[601] = 12'h777;
rom[602] = 12'h777;
rom[603] = 12'h777;
rom[604] = 12'h777;
rom[605] = 12'h777;
rom[606] = 12'h777;
rom[607] = 12'h777;
rom[608] = 12'h777;
rom[609] = 12'h777;
rom[610] = 12'h777;
rom[611] = 12'h777;
rom[612] = 12'h777;
rom[613] = 12'h777;
rom[614] = 12'h777;
rom[615] = 12'h777;
rom[616] = 12'h777;
rom[617] = 12'h777;
rom[618] = 12'h777;
rom[619] = 12'h777;
rom[620] = 12'h777;
rom[621] = 12'h777;
rom[622] = 12'h777;
rom[623] = 12'h777;
rom[624] = 12'h777;
  end
  endmodule


  module dash_rom (                       //тире
  input  wire    [13:0]     addr,
  output wire    [11:0]     word
);

  logic [11:0] rom [(46 * 26)];

  assign word = rom[addr];

  initial begin
rom[0] = 12'h000;
rom[1] = 12'h000;
rom[2] = 12'h000;
rom[3] = 12'h000;
rom[4] = 12'h000;
rom[5] = 12'h000;
rom[6] = 12'h000;
rom[7] = 12'h000;
rom[8] = 12'h000;
rom[9] = 12'h000;
rom[10] = 12'h000;
rom[11] = 12'h000;
rom[12] = 12'h000;
rom[13] = 12'h000;
rom[14] = 12'h000;
rom[15] = 12'h000;
rom[16] = 12'h000;
rom[17] = 12'h000;
rom[18] = 12'h000;
rom[19] = 12'h000;
rom[20] = 12'h000;
rom[21] = 12'h000;
rom[22] = 12'h000;
rom[23] = 12'h000;
rom[24] = 12'h000;
rom[25] = 12'h000;
rom[26] = 12'h000;
rom[27] = 12'h000;
rom[28] = 12'h000;
rom[29] = 12'h000;
rom[30] = 12'h000;
rom[31] = 12'h000;
rom[32] = 12'h000;
rom[33] = 12'h000;
rom[34] = 12'h000;
rom[35] = 12'h000;
rom[36] = 12'h000;
rom[37] = 12'h000;
rom[38] = 12'h000;
rom[39] = 12'h000;
rom[40] = 12'h000;
rom[41] = 12'h000;
rom[42] = 12'h000;
rom[43] = 12'h000;
rom[44] = 12'h000;
rom[45] = 12'h000;
rom[46] = 12'h000;
rom[47] = 12'h000;
rom[48] = 12'h000;
rom[49] = 12'h000;
rom[50] = 12'h000;
rom[51] = 12'h000;
rom[52] = 12'h000;
rom[53] = 12'h000;
rom[54] = 12'h000;
rom[55] = 12'h000;
rom[56] = 12'h000;
rom[57] = 12'h000;
rom[58] = 12'h007;
rom[59] = 12'h007;
rom[60] = 12'h000;
rom[61] = 12'h000;
rom[62] = 12'h007;
rom[63] = 12'h007;
rom[64] = 12'h000;
rom[65] = 12'h000;
rom[66] = 12'h007;
rom[67] = 12'h007;
rom[68] = 12'h000;
rom[69] = 12'h000;
rom[70] = 12'h007;
rom[71] = 12'h007;
rom[72] = 12'h000;
rom[73] = 12'h000;
rom[74] = 12'h000;
rom[75] = 12'h000;
rom[76] = 12'h000;
rom[77] = 12'h000;
rom[78] = 12'h000;
rom[79] = 12'h000;
rom[80] = 12'h000;
rom[81] = 12'h000;
rom[82] = 12'h000;
rom[83] = 12'h000;
rom[84] = 12'h007;
rom[85] = 12'h007;
rom[86] = 12'h000;
rom[87] = 12'h000;
rom[88] = 12'h007;
rom[89] = 12'h007;
rom[90] = 12'h000;
rom[91] = 12'h000;
rom[92] = 12'h007;
rom[93] = 12'h007;
rom[94] = 12'h000;
rom[95] = 12'h000;
rom[96] = 12'h007;
rom[97] = 12'h007;
rom[98] = 12'h000;
rom[99] = 12'h000;
rom[100] = 12'h000;
rom[101] = 12'h000;
rom[102] = 12'h000;
rom[103] = 12'h000;
rom[104] = 12'h000;
rom[105] = 12'h000;
rom[106] = 12'h007;
rom[107] = 12'h007;
rom[108] = 12'h000;
rom[109] = 12'h000;
rom[110] = 12'h000;
rom[111] = 12'h000;
rom[112] = 12'h007;
rom[113] = 12'h007;
rom[114] = 12'h000;
rom[115] = 12'h000;
rom[116] = 12'h007;
rom[117] = 12'h007;
rom[118] = 12'h000;
rom[119] = 12'h000;
rom[120] = 12'h007;
rom[121] = 12'h007;
rom[122] = 12'h000;
rom[123] = 12'h000;
rom[124] = 12'h000;
rom[125] = 12'h000;
rom[126] = 12'h007;
rom[127] = 12'h007;
rom[128] = 12'h000;
rom[129] = 12'h000;
rom[130] = 12'h000;
rom[131] = 12'h000;
rom[132] = 12'h007;
rom[133] = 12'h007;
rom[134] = 12'h000;
rom[135] = 12'h000;
rom[136] = 12'h000;
rom[137] = 12'h000;
rom[138] = 12'h007;
rom[139] = 12'h007;
rom[140] = 12'h000;
rom[141] = 12'h000;
rom[142] = 12'h007;
rom[143] = 12'h007;
rom[144] = 12'h000;
rom[145] = 12'h000;
rom[146] = 12'h007;
rom[147] = 12'h007;
rom[148] = 12'h000;
rom[149] = 12'h000;
rom[150] = 12'h000;
rom[151] = 12'h000;
rom[152] = 12'h007;
rom[153] = 12'h007;
rom[154] = 12'h000;
rom[155] = 12'h000;
rom[156] = 12'h000;
rom[157] = 12'h000;
rom[158] = 12'h000;
rom[159] = 12'h000;
rom[160] = 12'h007;
rom[161] = 12'h007;
rom[162] = 12'h000;
rom[163] = 12'h000;
rom[164] = 12'h000;
rom[165] = 12'h000;
rom[166] = 12'h007;
rom[167] = 12'h007;
rom[168] = 12'h000;
rom[169] = 12'h000;
rom[170] = 12'h007;
rom[171] = 12'h007;
rom[172] = 12'h000;
rom[173] = 12'h000;
rom[174] = 12'h000;
rom[175] = 12'h000;
rom[176] = 12'h007;
rom[177] = 12'h007;
rom[178] = 12'h000;
rom[179] = 12'h000;
rom[180] = 12'h000;
rom[181] = 12'h000;
rom[182] = 12'h000;
rom[183] = 12'h000;
rom[184] = 12'h000;
rom[185] = 12'h000;
rom[186] = 12'h007;
rom[187] = 12'h007;
rom[188] = 12'h000;
rom[189] = 12'h000;
rom[190] = 12'h000;
rom[191] = 12'h000;
rom[192] = 12'h007;
rom[193] = 12'h007;
rom[194] = 12'h000;
rom[195] = 12'h000;
rom[196] = 12'h007;
rom[197] = 12'h007;
rom[198] = 12'h000;
rom[199] = 12'h000;
rom[200] = 12'h000;
rom[201] = 12'h000;
rom[202] = 12'h007;
rom[203] = 12'h007;
rom[204] = 12'h000;
rom[205] = 12'h000;
rom[206] = 12'h000;
rom[207] = 12'h000;
rom[208] = 12'h000;
rom[209] = 12'h000;
rom[210] = 12'h007;
rom[211] = 12'h007;
rom[212] = 12'h000;
rom[213] = 12'h000;
rom[214] = 12'h007;
rom[215] = 12'h007;
rom[216] = 12'h000;
rom[217] = 12'h000;
rom[218] = 12'h000;
rom[219] = 12'h000;
rom[220] = 12'h000;
rom[221] = 12'h000;
rom[222] = 12'h000;
rom[223] = 12'h000;
rom[224] = 12'h000;
rom[225] = 12'h000;
rom[226] = 12'h007;
rom[227] = 12'h007;
rom[228] = 12'h000;
rom[229] = 12'h000;
rom[230] = 12'h007;
rom[231] = 12'h007;
rom[232] = 12'h000;
rom[233] = 12'h000;
rom[234] = 12'h000;
rom[235] = 12'h000;
rom[236] = 12'h007;
rom[237] = 12'h007;
rom[238] = 12'h000;
rom[239] = 12'h000;
rom[240] = 12'h007;
rom[241] = 12'h007;
rom[242] = 12'h000;
rom[243] = 12'h000;
rom[244] = 12'h000;
rom[245] = 12'h000;
rom[246] = 12'h000;
rom[247] = 12'h000;
rom[248] = 12'h000;
rom[249] = 12'h000;
rom[250] = 12'h000;
rom[251] = 12'h000;
rom[252] = 12'h007;
rom[253] = 12'h007;
rom[254] = 12'h000;
rom[255] = 12'h000;
rom[256] = 12'h007;
rom[257] = 12'h007;
rom[258] = 12'h000;
rom[259] = 12'h000;
rom[260] = 12'h000;
rom[261] = 12'h000;
rom[262] = 12'h000;
rom[263] = 12'h000;
rom[264] = 12'h007;
rom[265] = 12'h007;
rom[266] = 12'h000;
rom[267] = 12'h000;
rom[268] = 12'h000;
rom[269] = 12'h000;
rom[270] = 12'h000;
rom[271] = 12'h000;
rom[272] = 12'h000;
rom[273] = 12'h000;
rom[274] = 12'h000;
rom[275] = 12'h000;
rom[276] = 12'h000;
rom[277] = 12'h000;
rom[278] = 12'h000;
rom[279] = 12'h000;
rom[280] = 12'h007;
rom[281] = 12'h007;
rom[282] = 12'h000;
rom[283] = 12'h000;
rom[284] = 12'h000;
rom[285] = 12'h000;
rom[286] = 12'h000;
rom[287] = 12'h000;
rom[288] = 12'h000;
rom[289] = 12'h000;
rom[290] = 12'h007;
rom[291] = 12'h007;
rom[292] = 12'h000;
rom[293] = 12'h000;
rom[294] = 12'h000;
rom[295] = 12'h000;
rom[296] = 12'h000;
rom[297] = 12'h000;
rom[298] = 12'h000;
rom[299] = 12'h000;
rom[300] = 12'h000;
rom[301] = 12'h000;
rom[302] = 12'h000;
rom[303] = 12'h000;
rom[304] = 12'h000;
rom[305] = 12'h000;
rom[306] = 12'h007;
rom[307] = 12'h007;
rom[308] = 12'h000;
rom[309] = 12'h000;
rom[310] = 12'h000;
rom[311] = 12'h000;
rom[312] = 12'h000;
rom[313] = 12'h000;
rom[314] = 12'h007;
rom[315] = 12'h007;
rom[316] = 12'h000;
rom[317] = 12'h000;
rom[318] = 12'h007;
rom[319] = 12'h007;
rom[320] = 12'h000;
rom[321] = 12'h000;
rom[322] = 12'h000;
rom[323] = 12'h000;
rom[324] = 12'h000;
rom[325] = 12'h000;
rom[326] = 12'h000;
rom[327] = 12'h000;
rom[328] = 12'h000;
rom[329] = 12'h000;
rom[330] = 12'h007;
rom[331] = 12'h007;
rom[332] = 12'h000;
rom[333] = 12'h000;
rom[334] = 12'h007;
rom[335] = 12'h007;
rom[336] = 12'h000;
rom[337] = 12'h000;
rom[338] = 12'h000;
rom[339] = 12'h000;
rom[340] = 12'h007;
rom[341] = 12'h007;
rom[342] = 12'h000;
rom[343] = 12'h000;
rom[344] = 12'h007;
rom[345] = 12'h007;
rom[346] = 12'h000;
rom[347] = 12'h000;
rom[348] = 12'h000;
rom[349] = 12'h000;
rom[350] = 12'h000;
rom[351] = 12'h000;
rom[352] = 12'h000;
rom[353] = 12'h000;
rom[354] = 12'h000;
rom[355] = 12'h000;
rom[356] = 12'h007;
rom[357] = 12'h007;
rom[358] = 12'h000;
rom[359] = 12'h000;
rom[360] = 12'h007;
rom[361] = 12'h007;
rom[362] = 12'h000;
rom[363] = 12'h000;
rom[364] = 12'h000;
rom[365] = 12'h000;
rom[366] = 12'h000;
rom[367] = 12'h000;
rom[368] = 12'h007;
rom[369] = 12'h007;
rom[370] = 12'h000;
rom[371] = 12'h000;
rom[372] = 12'h000;
rom[373] = 12'h000;
rom[374] = 12'h000;
rom[375] = 12'h000;
rom[376] = 12'h000;
rom[377] = 12'h000;
rom[378] = 12'h000;
rom[379] = 12'h000;
rom[380] = 12'h000;
rom[381] = 12'h000;
rom[382] = 12'h000;
rom[383] = 12'h000;
rom[384] = 12'h007;
rom[385] = 12'h007;
rom[386] = 12'h000;
rom[387] = 12'h000;
rom[388] = 12'h000;
rom[389] = 12'h000;
rom[390] = 12'h000;
rom[391] = 12'h000;
rom[392] = 12'h000;
rom[393] = 12'h000;
rom[394] = 12'h007;
rom[395] = 12'h007;
rom[396] = 12'h000;
rom[397] = 12'h000;
rom[398] = 12'h000;
rom[399] = 12'h000;
rom[400] = 12'h000;
rom[401] = 12'h000;
rom[402] = 12'h000;
rom[403] = 12'h000;
rom[404] = 12'h000;
rom[405] = 12'h000;
rom[406] = 12'h000;
rom[407] = 12'h000;
rom[408] = 12'h000;
rom[409] = 12'h000;
rom[410] = 12'h007;
rom[411] = 12'h007;
rom[412] = 12'h000;
rom[413] = 12'h000;
rom[414] = 12'h000;
rom[415] = 12'h000;
rom[416] = 12'h000;
rom[417] = 12'h000;
rom[418] = 12'h007;
rom[419] = 12'h007;
rom[420] = 12'h000;
rom[421] = 12'h000;
rom[422] = 12'h007;
rom[423] = 12'h007;
rom[424] = 12'h000;
rom[425] = 12'h000;
rom[426] = 12'h000;
rom[427] = 12'h000;
rom[428] = 12'h000;
rom[429] = 12'h000;
rom[430] = 12'h000;
rom[431] = 12'h000;
rom[432] = 12'h000;
rom[433] = 12'h000;
rom[434] = 12'h007;
rom[435] = 12'h007;
rom[436] = 12'h000;
rom[437] = 12'h000;
rom[438] = 12'h007;
rom[439] = 12'h007;
rom[440] = 12'h000;
rom[441] = 12'h000;
rom[442] = 12'h000;
rom[443] = 12'h000;
rom[444] = 12'h007;
rom[445] = 12'h007;
rom[446] = 12'h000;
rom[447] = 12'h000;
rom[448] = 12'h007;
rom[449] = 12'h007;
rom[450] = 12'h000;
rom[451] = 12'h000;
rom[452] = 12'h000;
rom[453] = 12'h000;
rom[454] = 12'h000;
rom[455] = 12'h000;
rom[456] = 12'h000;
rom[457] = 12'h000;
rom[458] = 12'h000;
rom[459] = 12'h000;
rom[460] = 12'h007;
rom[461] = 12'h007;
rom[462] = 12'h000;
rom[463] = 12'h000;
rom[464] = 12'h007;
rom[465] = 12'h007;
rom[466] = 12'h000;
rom[467] = 12'h000;
rom[468] = 12'h000;
rom[469] = 12'h000;
rom[470] = 12'h000;
rom[471] = 12'h000;
rom[472] = 12'h007;
rom[473] = 12'h007;
rom[474] = 12'h000;
rom[475] = 12'h000;
rom[476] = 12'h000;
rom[477] = 12'h000;
rom[478] = 12'h000;
rom[479] = 12'h000;
rom[480] = 12'h000;
rom[481] = 12'h000;
rom[482] = 12'h000;
rom[483] = 12'h000;
rom[484] = 12'h000;
rom[485] = 12'h000;
rom[486] = 12'h000;
rom[487] = 12'h000;
rom[488] = 12'h007;
rom[489] = 12'h007;
rom[490] = 12'h000;
rom[491] = 12'h000;
rom[492] = 12'h000;
rom[493] = 12'h000;
rom[494] = 12'h000;
rom[495] = 12'h000;
rom[496] = 12'h000;
rom[497] = 12'h000;
rom[498] = 12'h007;
rom[499] = 12'h007;
rom[500] = 12'h000;
rom[501] = 12'h000;
rom[502] = 12'h000;
rom[503] = 12'h000;
rom[504] = 12'h000;
rom[505] = 12'h000;
rom[506] = 12'h000;
rom[507] = 12'h000;
rom[508] = 12'h000;
rom[509] = 12'h000;
rom[510] = 12'h000;
rom[511] = 12'h000;
rom[512] = 12'h000;
rom[513] = 12'h000;
rom[514] = 12'h007;
rom[515] = 12'h007;
rom[516] = 12'h000;
rom[517] = 12'h000;
rom[518] = 12'h000;
rom[519] = 12'h000;
rom[520] = 12'h000;
rom[521] = 12'h000;
rom[522] = 12'h007;
rom[523] = 12'h007;
rom[524] = 12'h000;
rom[525] = 12'h000;
rom[526] = 12'h00f;
rom[527] = 12'h00f;
rom[528] = 12'h00f;
rom[529] = 12'h00f;
rom[530] = 12'h00f;
rom[531] = 12'h00f;
rom[532] = 12'h00f;
rom[533] = 12'h00f;
rom[534] = 12'h00f;
rom[535] = 12'h00f;
rom[536] = 12'h00f;
rom[537] = 12'h00f;
rom[538] = 12'h00f;
rom[539] = 12'h00f;
rom[540] = 12'h000;
rom[541] = 12'h000;
rom[542] = 12'h007;
rom[543] = 12'h007;
rom[544] = 12'h000;
rom[545] = 12'h000;
rom[546] = 12'h000;
rom[547] = 12'h000;
rom[548] = 12'h007;
rom[549] = 12'h007;
rom[550] = 12'h000;
rom[551] = 12'h000;
rom[552] = 12'h00f;
rom[553] = 12'h00f;
rom[554] = 12'h00f;
rom[555] = 12'h00f;
rom[556] = 12'h00f;
rom[557] = 12'h00f;
rom[558] = 12'h00f;
rom[559] = 12'h00f;
rom[560] = 12'h00f;
rom[561] = 12'h00f;
rom[562] = 12'h00f;
rom[563] = 12'h00f;
rom[564] = 12'h00f;
rom[565] = 12'h00f;
rom[566] = 12'h000;
rom[567] = 12'h000;
rom[568] = 12'h007;
rom[569] = 12'h007;
rom[570] = 12'h000;
rom[571] = 12'h000;
rom[572] = 12'h000;
rom[573] = 12'h000;
rom[574] = 12'h000;
rom[575] = 12'h000;
rom[576] = 12'h00f;
rom[577] = 12'h00f;
rom[578] = 12'h00f;
rom[579] = 12'h00f;
rom[580] = 12'h00f;
rom[581] = 12'h00f;
rom[582] = 12'h00f;
rom[583] = 12'h00f;
rom[584] = 12'h00f;
rom[585] = 12'h00f;
rom[586] = 12'h00f;
rom[587] = 12'h00f;
rom[588] = 12'h00f;
rom[589] = 12'h00f;
rom[590] = 12'h00f;
rom[591] = 12'h00f;
rom[592] = 12'h00f;
rom[593] = 12'h00f;
rom[594] = 12'h000;
rom[595] = 12'h000;
rom[596] = 12'h000;
rom[597] = 12'h000;
rom[598] = 12'h000;
rom[599] = 12'h000;
rom[600] = 12'h000;
rom[601] = 12'h000;
rom[602] = 12'h00f;
rom[603] = 12'h00f;
rom[604] = 12'h00f;
rom[605] = 12'h00f;
rom[606] = 12'h00f;
rom[607] = 12'h00f;
rom[608] = 12'h00f;
rom[609] = 12'h00f;
rom[610] = 12'h00f;
rom[611] = 12'h00f;
rom[612] = 12'h00f;
rom[613] = 12'h00f;
rom[614] = 12'h00f;
rom[615] = 12'h00f;
rom[616] = 12'h00f;
rom[617] = 12'h00f;
rom[618] = 12'h00f;
rom[619] = 12'h00f;
rom[620] = 12'h000;
rom[621] = 12'h000;
rom[622] = 12'h000;
rom[623] = 12'h000;
rom[624] = 12'h000;
rom[625] = 12'h000;
rom[626] = 12'h007;
rom[627] = 12'h007;
rom[628] = 12'h000;
rom[629] = 12'h000;
rom[630] = 12'h00f;
rom[631] = 12'h00f;
rom[632] = 12'h00f;
rom[633] = 12'h00f;
rom[634] = 12'h00f;
rom[635] = 12'h00f;
rom[636] = 12'h00f;
rom[637] = 12'h00f;
rom[638] = 12'h00f;
rom[639] = 12'h00f;
rom[640] = 12'h00f;
rom[641] = 12'h00f;
rom[642] = 12'h00f;
rom[643] = 12'h00f;
rom[644] = 12'h000;
rom[645] = 12'h000;
rom[646] = 12'h007;
rom[647] = 12'h007;
rom[648] = 12'h000;
rom[649] = 12'h000;
rom[650] = 12'h000;
rom[651] = 12'h000;
rom[652] = 12'h007;
rom[653] = 12'h007;
rom[654] = 12'h000;
rom[655] = 12'h000;
rom[656] = 12'h00f;
rom[657] = 12'h00f;
rom[658] = 12'h00f;
rom[659] = 12'h00f;
rom[660] = 12'h00f;
rom[661] = 12'h00f;
rom[662] = 12'h00f;
rom[663] = 12'h00f;
rom[664] = 12'h00f;
rom[665] = 12'h00f;
rom[666] = 12'h00f;
rom[667] = 12'h00f;
rom[668] = 12'h00f;
rom[669] = 12'h00f;
rom[670] = 12'h000;
rom[671] = 12'h000;
rom[672] = 12'h007;
rom[673] = 12'h007;
rom[674] = 12'h000;
rom[675] = 12'h000;
rom[676] = 12'h000;
rom[677] = 12'h000;
rom[678] = 12'h000;
rom[679] = 12'h000;
rom[680] = 12'h007;
rom[681] = 12'h007;
rom[682] = 12'h000;
rom[683] = 12'h000;
rom[684] = 12'h000;
rom[685] = 12'h000;
rom[686] = 12'h000;
rom[687] = 12'h000;
rom[688] = 12'h000;
rom[689] = 12'h000;
rom[690] = 12'h000;
rom[691] = 12'h000;
rom[692] = 12'h000;
rom[693] = 12'h000;
rom[694] = 12'h000;
rom[695] = 12'h000;
rom[696] = 12'h007;
rom[697] = 12'h007;
rom[698] = 12'h000;
rom[699] = 12'h000;
rom[700] = 12'h000;
rom[701] = 12'h000;
rom[702] = 12'h000;
rom[703] = 12'h000;
rom[704] = 12'h000;
rom[705] = 12'h000;
rom[706] = 12'h007;
rom[707] = 12'h007;
rom[708] = 12'h000;
rom[709] = 12'h000;
rom[710] = 12'h000;
rom[711] = 12'h000;
rom[712] = 12'h000;
rom[713] = 12'h000;
rom[714] = 12'h000;
rom[715] = 12'h000;
rom[716] = 12'h000;
rom[717] = 12'h000;
rom[718] = 12'h000;
rom[719] = 12'h000;
rom[720] = 12'h000;
rom[721] = 12'h000;
rom[722] = 12'h007;
rom[723] = 12'h007;
rom[724] = 12'h000;
rom[725] = 12'h000;
rom[726] = 12'h000;
rom[727] = 12'h000;
rom[728] = 12'h000;
rom[729] = 12'h000;
rom[730] = 12'h007;
rom[731] = 12'h007;
rom[732] = 12'h000;
rom[733] = 12'h000;
rom[734] = 12'h007;
rom[735] = 12'h007;
rom[736] = 12'h000;
rom[737] = 12'h000;
rom[738] = 12'h000;
rom[739] = 12'h000;
rom[740] = 12'h000;
rom[741] = 12'h000;
rom[742] = 12'h000;
rom[743] = 12'h000;
rom[744] = 12'h000;
rom[745] = 12'h000;
rom[746] = 12'h007;
rom[747] = 12'h007;
rom[748] = 12'h000;
rom[749] = 12'h000;
rom[750] = 12'h007;
rom[751] = 12'h007;
rom[752] = 12'h000;
rom[753] = 12'h000;
rom[754] = 12'h000;
rom[755] = 12'h000;
rom[756] = 12'h007;
rom[757] = 12'h007;
rom[758] = 12'h000;
rom[759] = 12'h000;
rom[760] = 12'h007;
rom[761] = 12'h007;
rom[762] = 12'h000;
rom[763] = 12'h000;
rom[764] = 12'h000;
rom[765] = 12'h000;
rom[766] = 12'h000;
rom[767] = 12'h000;
rom[768] = 12'h000;
rom[769] = 12'h000;
rom[770] = 12'h000;
rom[771] = 12'h000;
rom[772] = 12'h007;
rom[773] = 12'h007;
rom[774] = 12'h000;
rom[775] = 12'h000;
rom[776] = 12'h007;
rom[777] = 12'h007;
rom[778] = 12'h000;
rom[779] = 12'h000;
rom[780] = 12'h000;
rom[781] = 12'h000;
rom[782] = 12'h000;
rom[783] = 12'h000;
rom[784] = 12'h007;
rom[785] = 12'h007;
rom[786] = 12'h000;
rom[787] = 12'h000;
rom[788] = 12'h000;
rom[789] = 12'h000;
rom[790] = 12'h000;
rom[791] = 12'h000;
rom[792] = 12'h000;
rom[793] = 12'h000;
rom[794] = 12'h000;
rom[795] = 12'h000;
rom[796] = 12'h000;
rom[797] = 12'h000;
rom[798] = 12'h000;
rom[799] = 12'h000;
rom[800] = 12'h007;
rom[801] = 12'h007;
rom[802] = 12'h000;
rom[803] = 12'h000;
rom[804] = 12'h000;
rom[805] = 12'h000;
rom[806] = 12'h000;
rom[807] = 12'h000;
rom[808] = 12'h000;
rom[809] = 12'h000;
rom[810] = 12'h007;
rom[811] = 12'h007;
rom[812] = 12'h000;
rom[813] = 12'h000;
rom[814] = 12'h000;
rom[815] = 12'h000;
rom[816] = 12'h000;
rom[817] = 12'h000;
rom[818] = 12'h000;
rom[819] = 12'h000;
rom[820] = 12'h000;
rom[821] = 12'h000;
rom[822] = 12'h000;
rom[823] = 12'h000;
rom[824] = 12'h000;
rom[825] = 12'h000;
rom[826] = 12'h007;
rom[827] = 12'h007;
rom[828] = 12'h000;
rom[829] = 12'h000;
rom[830] = 12'h000;
rom[831] = 12'h000;
rom[832] = 12'h000;
rom[833] = 12'h000;
rom[834] = 12'h007;
rom[835] = 12'h007;
rom[836] = 12'h000;
rom[837] = 12'h000;
rom[838] = 12'h007;
rom[839] = 12'h007;
rom[840] = 12'h000;
rom[841] = 12'h000;
rom[842] = 12'h000;
rom[843] = 12'h000;
rom[844] = 12'h000;
rom[845] = 12'h000;
rom[846] = 12'h000;
rom[847] = 12'h000;
rom[848] = 12'h000;
rom[849] = 12'h000;
rom[850] = 12'h007;
rom[851] = 12'h007;
rom[852] = 12'h000;
rom[853] = 12'h000;
rom[854] = 12'h007;
rom[855] = 12'h007;
rom[856] = 12'h000;
rom[857] = 12'h000;
rom[858] = 12'h000;
rom[859] = 12'h000;
rom[860] = 12'h007;
rom[861] = 12'h007;
rom[862] = 12'h000;
rom[863] = 12'h000;
rom[864] = 12'h007;
rom[865] = 12'h007;
rom[866] = 12'h000;
rom[867] = 12'h000;
rom[868] = 12'h000;
rom[869] = 12'h000;
rom[870] = 12'h000;
rom[871] = 12'h000;
rom[872] = 12'h000;
rom[873] = 12'h000;
rom[874] = 12'h000;
rom[875] = 12'h000;
rom[876] = 12'h007;
rom[877] = 12'h007;
rom[878] = 12'h000;
rom[879] = 12'h000;
rom[880] = 12'h007;
rom[881] = 12'h007;
rom[882] = 12'h000;
rom[883] = 12'h000;
rom[884] = 12'h000;
rom[885] = 12'h000;
rom[886] = 12'h000;
rom[887] = 12'h000;
rom[888] = 12'h007;
rom[889] = 12'h007;
rom[890] = 12'h000;
rom[891] = 12'h000;
rom[892] = 12'h000;
rom[893] = 12'h000;
rom[894] = 12'h000;
rom[895] = 12'h000;
rom[896] = 12'h000;
rom[897] = 12'h000;
rom[898] = 12'h000;
rom[899] = 12'h000;
rom[900] = 12'h000;
rom[901] = 12'h000;
rom[902] = 12'h000;
rom[903] = 12'h000;
rom[904] = 12'h007;
rom[905] = 12'h007;
rom[906] = 12'h000;
rom[907] = 12'h000;
rom[908] = 12'h000;
rom[909] = 12'h000;
rom[910] = 12'h000;
rom[911] = 12'h000;
rom[912] = 12'h000;
rom[913] = 12'h000;
rom[914] = 12'h007;
rom[915] = 12'h007;
rom[916] = 12'h000;
rom[917] = 12'h000;
rom[918] = 12'h000;
rom[919] = 12'h000;
rom[920] = 12'h000;
rom[921] = 12'h000;
rom[922] = 12'h000;
rom[923] = 12'h000;
rom[924] = 12'h000;
rom[925] = 12'h000;
rom[926] = 12'h000;
rom[927] = 12'h000;
rom[928] = 12'h000;
rom[929] = 12'h000;
rom[930] = 12'h007;
rom[931] = 12'h007;
rom[932] = 12'h000;
rom[933] = 12'h000;
rom[934] = 12'h000;
rom[935] = 12'h000;
rom[936] = 12'h000;
rom[937] = 12'h000;
rom[938] = 12'h007;
rom[939] = 12'h007;
rom[940] = 12'h000;
rom[941] = 12'h000;
rom[942] = 12'h007;
rom[943] = 12'h007;
rom[944] = 12'h000;
rom[945] = 12'h000;
rom[946] = 12'h000;
rom[947] = 12'h000;
rom[948] = 12'h000;
rom[949] = 12'h000;
rom[950] = 12'h000;
rom[951] = 12'h000;
rom[952] = 12'h000;
rom[953] = 12'h000;
rom[954] = 12'h007;
rom[955] = 12'h007;
rom[956] = 12'h000;
rom[957] = 12'h000;
rom[958] = 12'h007;
rom[959] = 12'h007;
rom[960] = 12'h000;
rom[961] = 12'h000;
rom[962] = 12'h000;
rom[963] = 12'h000;
rom[964] = 12'h007;
rom[965] = 12'h007;
rom[966] = 12'h000;
rom[967] = 12'h000;
rom[968] = 12'h007;
rom[969] = 12'h007;
rom[970] = 12'h000;
rom[971] = 12'h000;
rom[972] = 12'h000;
rom[973] = 12'h000;
rom[974] = 12'h000;
rom[975] = 12'h000;
rom[976] = 12'h000;
rom[977] = 12'h000;
rom[978] = 12'h000;
rom[979] = 12'h000;
rom[980] = 12'h007;
rom[981] = 12'h007;
rom[982] = 12'h000;
rom[983] = 12'h000;
rom[984] = 12'h007;
rom[985] = 12'h007;
rom[986] = 12'h000;
rom[987] = 12'h000;
rom[988] = 12'h000;
rom[989] = 12'h000;
rom[990] = 12'h000;
rom[991] = 12'h000;
rom[992] = 12'h007;
rom[993] = 12'h007;
rom[994] = 12'h000;
rom[995] = 12'h000;
rom[996] = 12'h000;
rom[997] = 12'h000;
rom[998] = 12'h007;
rom[999] = 12'h007;
rom[1000] = 12'h000;
rom[1001] = 12'h000;
rom[1002] = 12'h007;
rom[1003] = 12'h007;
rom[1004] = 12'h000;
rom[1005] = 12'h000;
rom[1006] = 12'h000;
rom[1007] = 12'h000;
rom[1008] = 12'h007;
rom[1009] = 12'h007;
rom[1010] = 12'h000;
rom[1011] = 12'h000;
rom[1012] = 12'h000;
rom[1013] = 12'h000;
rom[1014] = 12'h000;
rom[1015] = 12'h000;
rom[1016] = 12'h000;
rom[1017] = 12'h000;
rom[1018] = 12'h007;
rom[1019] = 12'h007;
rom[1020] = 12'h000;
rom[1021] = 12'h000;
rom[1022] = 12'h000;
rom[1023] = 12'h000;
rom[1024] = 12'h007;
rom[1025] = 12'h007;
rom[1026] = 12'h000;
rom[1027] = 12'h000;
rom[1028] = 12'h007;
rom[1029] = 12'h007;
rom[1030] = 12'h000;
rom[1031] = 12'h000;
rom[1032] = 12'h000;
rom[1033] = 12'h000;
rom[1034] = 12'h007;
rom[1035] = 12'h007;
rom[1036] = 12'h000;
rom[1037] = 12'h000;
rom[1038] = 12'h000;
rom[1039] = 12'h000;
rom[1040] = 12'h000;
rom[1041] = 12'h000;
rom[1042] = 12'h007;
rom[1043] = 12'h007;
rom[1044] = 12'h000;
rom[1045] = 12'h000;
rom[1046] = 12'h000;
rom[1047] = 12'h000;
rom[1048] = 12'h007;
rom[1049] = 12'h007;
rom[1050] = 12'h000;
rom[1051] = 12'h000;
rom[1052] = 12'h007;
rom[1053] = 12'h007;
rom[1054] = 12'h000;
rom[1055] = 12'h000;
rom[1056] = 12'h007;
rom[1057] = 12'h007;
rom[1058] = 12'h000;
rom[1059] = 12'h000;
rom[1060] = 12'h000;
rom[1061] = 12'h000;
rom[1062] = 12'h007;
rom[1063] = 12'h007;
rom[1064] = 12'h000;
rom[1065] = 12'h000;
rom[1066] = 12'h000;
rom[1067] = 12'h000;
rom[1068] = 12'h007;
rom[1069] = 12'h007;
rom[1070] = 12'h000;
rom[1071] = 12'h000;
rom[1072] = 12'h000;
rom[1073] = 12'h000;
rom[1074] = 12'h007;
rom[1075] = 12'h007;
rom[1076] = 12'h000;
rom[1077] = 12'h000;
rom[1078] = 12'h007;
rom[1079] = 12'h007;
rom[1080] = 12'h000;
rom[1081] = 12'h000;
rom[1082] = 12'h007;
rom[1083] = 12'h007;
rom[1084] = 12'h000;
rom[1085] = 12'h000;
rom[1086] = 12'h000;
rom[1087] = 12'h000;
rom[1088] = 12'h007;
rom[1089] = 12'h007;
rom[1090] = 12'h000;
rom[1091] = 12'h000;
rom[1092] = 12'h000;
rom[1093] = 12'h000;
rom[1094] = 12'h000;
rom[1095] = 12'h000;
rom[1096] = 12'h000;
rom[1097] = 12'h000;
rom[1098] = 12'h007;
rom[1099] = 12'h007;
rom[1100] = 12'h000;
rom[1101] = 12'h000;
rom[1102] = 12'h007;
rom[1103] = 12'h007;
rom[1104] = 12'h000;
rom[1105] = 12'h000;
rom[1106] = 12'h007;
rom[1107] = 12'h007;
rom[1108] = 12'h000;
rom[1109] = 12'h000;
rom[1110] = 12'h007;
rom[1111] = 12'h007;
rom[1112] = 12'h000;
rom[1113] = 12'h000;
rom[1114] = 12'h000;
rom[1115] = 12'h000;
rom[1116] = 12'h000;
rom[1117] = 12'h000;
rom[1118] = 12'h000;
rom[1119] = 12'h000;
rom[1120] = 12'h000;
rom[1121] = 12'h000;
rom[1122] = 12'h000;
rom[1123] = 12'h000;
rom[1124] = 12'h007;
rom[1125] = 12'h007;
rom[1126] = 12'h000;
rom[1127] = 12'h000;
rom[1128] = 12'h007;
rom[1129] = 12'h007;
rom[1130] = 12'h000;
rom[1131] = 12'h000;
rom[1132] = 12'h007;
rom[1133] = 12'h007;
rom[1134] = 12'h000;
rom[1135] = 12'h000;
rom[1136] = 12'h007;
rom[1137] = 12'h007;
rom[1138] = 12'h000;
rom[1139] = 12'h000;
rom[1140] = 12'h000;
rom[1141] = 12'h000;
rom[1142] = 12'h000;
rom[1143] = 12'h000;
rom[1144] = 12'h000;
rom[1145] = 12'h000;
rom[1146] = 12'h000;
rom[1147] = 12'h000;
rom[1148] = 12'h000;
rom[1149] = 12'h000;
rom[1150] = 12'h000;
rom[1151] = 12'h000;
rom[1152] = 12'h000;
rom[1153] = 12'h000;
rom[1154] = 12'h000;
rom[1155] = 12'h000;
rom[1156] = 12'h000;
rom[1157] = 12'h000;
rom[1158] = 12'h000;
rom[1159] = 12'h000;
rom[1160] = 12'h000;
rom[1161] = 12'h000;
rom[1162] = 12'h000;
rom[1163] = 12'h000;
rom[1164] = 12'h000;
rom[1165] = 12'h000;
rom[1166] = 12'h000;
rom[1167] = 12'h000;
rom[1168] = 12'h000;
rom[1169] = 12'h000;
rom[1170] = 12'h000;
rom[1171] = 12'h000;
rom[1172] = 12'h000;
rom[1173] = 12'h000;
rom[1174] = 12'h000;
rom[1175] = 12'h000;
rom[1176] = 12'h000;
rom[1177] = 12'h000;
rom[1178] = 12'h000;
rom[1179] = 12'h000;
rom[1180] = 12'h000;
rom[1181] = 12'h000;
rom[1182] = 12'h000;
rom[1183] = 12'h000;
rom[1184] = 12'h000;
rom[1185] = 12'h000;
rom[1186] = 12'h000;
rom[1187] = 12'h000;
rom[1188] = 12'h000;
rom[1189] = 12'h000;
rom[1190] = 12'h000;
rom[1191] = 12'h000;
rom[1192] = 12'h000;
rom[1193] = 12'h000;
rom[1194] = 12'h000;
rom[1195] = 12'h000;
  end
  endmodule

    module zero_rom (                       //ноль
  input  wire    [13:0]     addr,
  output wire    [11:0]     word
);

  logic [11:0] rom [(46 * 26)];

  assign word = rom[addr];

  initial begin
rom[0] = 12'h000;
rom[1] = 12'h000;
rom[2] = 12'h000;
rom[3] = 12'h000;
rom[4] = 12'h000;
rom[5] = 12'h000;
rom[6] = 12'h000;
rom[7] = 12'h000;
rom[8] = 12'h000;
rom[9] = 12'h000;
rom[10] = 12'h000;
rom[11] = 12'h000;
rom[12] = 12'h000;
rom[13] = 12'h000;
rom[14] = 12'h000;
rom[15] = 12'h000;
rom[16] = 12'h000;
rom[17] = 12'h000;
rom[18] = 12'h000;
rom[19] = 12'h000;
rom[20] = 12'h000;
rom[21] = 12'h000;
rom[22] = 12'h000;
rom[23] = 12'h000;
rom[24] = 12'h000;
rom[25] = 12'h000;
rom[26] = 12'h000;
rom[27] = 12'h000;
rom[28] = 12'h000;
rom[29] = 12'h000;
rom[30] = 12'h000;
rom[31] = 12'h000;
rom[32] = 12'h000;
rom[33] = 12'h000;
rom[34] = 12'h000;
rom[35] = 12'h000;
rom[36] = 12'h000;
rom[37] = 12'h000;
rom[38] = 12'h000;
rom[39] = 12'h000;
rom[40] = 12'h000;
rom[41] = 12'h000;
rom[42] = 12'h000;
rom[43] = 12'h000;
rom[44] = 12'h000;
rom[45] = 12'h000;
rom[46] = 12'h000;
rom[47] = 12'h000;
rom[48] = 12'h000;
rom[49] = 12'h000;
rom[50] = 12'h000;
rom[51] = 12'h000;
rom[52] = 12'h000;
rom[53] = 12'h000;
rom[54] = 12'h000;
rom[55] = 12'h000;
rom[56] = 12'h00f;
rom[57] = 12'h00f;
rom[58] = 12'h00f;
rom[59] = 12'h00f;
rom[60] = 12'h00f;
rom[61] = 12'h00f;
rom[62] = 12'h00f;
rom[63] = 12'h00f;
rom[64] = 12'h00f;
rom[65] = 12'h00f;
rom[66] = 12'h00f;
rom[67] = 12'h00f;
rom[68] = 12'h00f;
rom[69] = 12'h00f;
rom[70] = 12'h00f;
rom[71] = 12'h00f;
rom[72] = 12'h00f;
rom[73] = 12'h00f;
rom[74] = 12'h000;
rom[75] = 12'h000;
rom[76] = 12'h000;
rom[77] = 12'h000;
rom[78] = 12'h000;
rom[79] = 12'h000;
rom[80] = 12'h000;
rom[81] = 12'h000;
rom[82] = 12'h00f;
rom[83] = 12'h00f;
rom[84] = 12'h00f;
rom[85] = 12'h00f;
rom[86] = 12'h00f;
rom[87] = 12'h00f;
rom[88] = 12'h00f;
rom[89] = 12'h00f;
rom[90] = 12'h00f;
rom[91] = 12'h00f;
rom[92] = 12'h00f;
rom[93] = 12'h00f;
rom[94] = 12'h00f;
rom[95] = 12'h00f;
rom[96] = 12'h00f;
rom[97] = 12'h00f;
rom[98] = 12'h00f;
rom[99] = 12'h00f;
rom[100] = 12'h000;
rom[101] = 12'h000;
rom[102] = 12'h000;
rom[103] = 12'h000;
rom[104] = 12'h000;
rom[105] = 12'h000;
rom[106] = 12'h00f;
rom[107] = 12'h00f;
rom[108] = 12'h000;
rom[109] = 12'h000;
rom[110] = 12'h00f;
rom[111] = 12'h00f;
rom[112] = 12'h00f;
rom[113] = 12'h00f;
rom[114] = 12'h00f;
rom[115] = 12'h00f;
rom[116] = 12'h00f;
rom[117] = 12'h00f;
rom[118] = 12'h00f;
rom[119] = 12'h00f;
rom[120] = 12'h00f;
rom[121] = 12'h00f;
rom[122] = 12'h00f;
rom[123] = 12'h00f;
rom[124] = 12'h000;
rom[125] = 12'h000;
rom[126] = 12'h00f;
rom[127] = 12'h00f;
rom[128] = 12'h000;
rom[129] = 12'h000;
rom[130] = 12'h000;
rom[131] = 12'h000;
rom[132] = 12'h00f;
rom[133] = 12'h00f;
rom[134] = 12'h000;
rom[135] = 12'h000;
rom[136] = 12'h00f;
rom[137] = 12'h00f;
rom[138] = 12'h00f;
rom[139] = 12'h00f;
rom[140] = 12'h00f;
rom[141] = 12'h00f;
rom[142] = 12'h00f;
rom[143] = 12'h00f;
rom[144] = 12'h00f;
rom[145] = 12'h00f;
rom[146] = 12'h00f;
rom[147] = 12'h00f;
rom[148] = 12'h00f;
rom[149] = 12'h00f;
rom[150] = 12'h000;
rom[151] = 12'h000;
rom[152] = 12'h00f;
rom[153] = 12'h00f;
rom[154] = 12'h000;
rom[155] = 12'h000;
rom[156] = 12'h000;
rom[157] = 12'h000;
rom[158] = 12'h00f;
rom[159] = 12'h00f;
rom[160] = 12'h00f;
rom[161] = 12'h00f;
rom[162] = 12'h000;
rom[163] = 12'h000;
rom[164] = 12'h00f;
rom[165] = 12'h00f;
rom[166] = 12'h00f;
rom[167] = 12'h00f;
rom[168] = 12'h00f;
rom[169] = 12'h00f;
rom[170] = 12'h00f;
rom[171] = 12'h00f;
rom[172] = 12'h00f;
rom[173] = 12'h00f;
rom[174] = 12'h000;
rom[175] = 12'h000;
rom[176] = 12'h00f;
rom[177] = 12'h00f;
rom[178] = 12'h00f;
rom[179] = 12'h00f;
rom[180] = 12'h000;
rom[181] = 12'h000;
rom[182] = 12'h000;
rom[183] = 12'h000;
rom[184] = 12'h00f;
rom[185] = 12'h00f;
rom[186] = 12'h00f;
rom[187] = 12'h00f;
rom[188] = 12'h000;
rom[189] = 12'h000;
rom[190] = 12'h00f;
rom[191] = 12'h00f;
rom[192] = 12'h00f;
rom[193] = 12'h00f;
rom[194] = 12'h00f;
rom[195] = 12'h00f;
rom[196] = 12'h00f;
rom[197] = 12'h00f;
rom[198] = 12'h00f;
rom[199] = 12'h00f;
rom[200] = 12'h000;
rom[201] = 12'h000;
rom[202] = 12'h00f;
rom[203] = 12'h00f;
rom[204] = 12'h00f;
rom[205] = 12'h00f;
rom[206] = 12'h000;
rom[207] = 12'h000;
rom[208] = 12'h000;
rom[209] = 12'h000;
rom[210] = 12'h00f;
rom[211] = 12'h00f;
rom[212] = 12'h00f;
rom[213] = 12'h00f;
rom[214] = 12'h00f;
rom[215] = 12'h00f;
rom[216] = 12'h000;
rom[217] = 12'h000;
rom[218] = 12'h000;
rom[219] = 12'h000;
rom[220] = 12'h000;
rom[221] = 12'h000;
rom[222] = 12'h000;
rom[223] = 12'h000;
rom[224] = 12'h000;
rom[225] = 12'h000;
rom[226] = 12'h00f;
rom[227] = 12'h00f;
rom[228] = 12'h00f;
rom[229] = 12'h00f;
rom[230] = 12'h00f;
rom[231] = 12'h00f;
rom[232] = 12'h000;
rom[233] = 12'h000;
rom[234] = 12'h000;
rom[235] = 12'h000;
rom[236] = 12'h00f;
rom[237] = 12'h00f;
rom[238] = 12'h00f;
rom[239] = 12'h00f;
rom[240] = 12'h00f;
rom[241] = 12'h00f;
rom[242] = 12'h000;
rom[243] = 12'h000;
rom[244] = 12'h000;
rom[245] = 12'h000;
rom[246] = 12'h000;
rom[247] = 12'h000;
rom[248] = 12'h000;
rom[249] = 12'h000;
rom[250] = 12'h000;
rom[251] = 12'h000;
rom[252] = 12'h00f;
rom[253] = 12'h00f;
rom[254] = 12'h00f;
rom[255] = 12'h00f;
rom[256] = 12'h00f;
rom[257] = 12'h00f;
rom[258] = 12'h000;
rom[259] = 12'h000;
rom[260] = 12'h000;
rom[261] = 12'h000;
rom[262] = 12'h00f;
rom[263] = 12'h00f;
rom[264] = 12'h00f;
rom[265] = 12'h00f;
rom[266] = 12'h00f;
rom[267] = 12'h00f;
rom[268] = 12'h000;
rom[269] = 12'h000;
rom[270] = 12'h000;
rom[271] = 12'h000;
rom[272] = 12'h000;
rom[273] = 12'h000;
rom[274] = 12'h000;
rom[275] = 12'h000;
rom[276] = 12'h000;
rom[277] = 12'h000;
rom[278] = 12'h00f;
rom[279] = 12'h00f;
rom[280] = 12'h00f;
rom[281] = 12'h00f;
rom[282] = 12'h00f;
rom[283] = 12'h00f;
rom[284] = 12'h000;
rom[285] = 12'h000;
rom[286] = 12'h000;
rom[287] = 12'h000;
rom[288] = 12'h00f;
rom[289] = 12'h00f;
rom[290] = 12'h00f;
rom[291] = 12'h00f;
rom[292] = 12'h00f;
rom[293] = 12'h00f;
rom[294] = 12'h000;
rom[295] = 12'h000;
rom[296] = 12'h000;
rom[297] = 12'h000;
rom[298] = 12'h000;
rom[299] = 12'h000;
rom[300] = 12'h000;
rom[301] = 12'h000;
rom[302] = 12'h000;
rom[303] = 12'h000;
rom[304] = 12'h00f;
rom[305] = 12'h00f;
rom[306] = 12'h00f;
rom[307] = 12'h00f;
rom[308] = 12'h00f;
rom[309] = 12'h00f;
rom[310] = 12'h000;
rom[311] = 12'h000;
rom[312] = 12'h000;
rom[313] = 12'h000;
rom[314] = 12'h00f;
rom[315] = 12'h00f;
rom[316] = 12'h00f;
rom[317] = 12'h00f;
rom[318] = 12'h00f;
rom[319] = 12'h00f;
rom[320] = 12'h000;
rom[321] = 12'h000;
rom[322] = 12'h000;
rom[323] = 12'h000;
rom[324] = 12'h000;
rom[325] = 12'h000;
rom[326] = 12'h000;
rom[327] = 12'h000;
rom[328] = 12'h000;
rom[329] = 12'h000;
rom[330] = 12'h00f;
rom[331] = 12'h00f;
rom[332] = 12'h00f;
rom[333] = 12'h00f;
rom[334] = 12'h00f;
rom[335] = 12'h00f;
rom[336] = 12'h000;
rom[337] = 12'h000;
rom[338] = 12'h000;
rom[339] = 12'h000;
rom[340] = 12'h00f;
rom[341] = 12'h00f;
rom[342] = 12'h00f;
rom[343] = 12'h00f;
rom[344] = 12'h00f;
rom[345] = 12'h00f;
rom[346] = 12'h000;
rom[347] = 12'h000;
rom[348] = 12'h000;
rom[349] = 12'h000;
rom[350] = 12'h000;
rom[351] = 12'h000;
rom[352] = 12'h000;
rom[353] = 12'h000;
rom[354] = 12'h000;
rom[355] = 12'h000;
rom[356] = 12'h00f;
rom[357] = 12'h00f;
rom[358] = 12'h00f;
rom[359] = 12'h00f;
rom[360] = 12'h00f;
rom[361] = 12'h00f;
rom[362] = 12'h000;
rom[363] = 12'h000;
rom[364] = 12'h000;
rom[365] = 12'h000;
rom[366] = 12'h00f;
rom[367] = 12'h00f;
rom[368] = 12'h00f;
rom[369] = 12'h00f;
rom[370] = 12'h00f;
rom[371] = 12'h00f;
rom[372] = 12'h000;
rom[373] = 12'h000;
rom[374] = 12'h000;
rom[375] = 12'h000;
rom[376] = 12'h000;
rom[377] = 12'h000;
rom[378] = 12'h000;
rom[379] = 12'h000;
rom[380] = 12'h000;
rom[381] = 12'h000;
rom[382] = 12'h00f;
rom[383] = 12'h00f;
rom[384] = 12'h00f;
rom[385] = 12'h00f;
rom[386] = 12'h00f;
rom[387] = 12'h00f;
rom[388] = 12'h000;
rom[389] = 12'h000;
rom[390] = 12'h000;
rom[391] = 12'h000;
rom[392] = 12'h00f;
rom[393] = 12'h00f;
rom[394] = 12'h00f;
rom[395] = 12'h00f;
rom[396] = 12'h00f;
rom[397] = 12'h00f;
rom[398] = 12'h000;
rom[399] = 12'h000;
rom[400] = 12'h000;
rom[401] = 12'h000;
rom[402] = 12'h000;
rom[403] = 12'h000;
rom[404] = 12'h000;
rom[405] = 12'h000;
rom[406] = 12'h000;
rom[407] = 12'h000;
rom[408] = 12'h00f;
rom[409] = 12'h00f;
rom[410] = 12'h00f;
rom[411] = 12'h00f;
rom[412] = 12'h00f;
rom[413] = 12'h00f;
rom[414] = 12'h000;
rom[415] = 12'h000;
rom[416] = 12'h000;
rom[417] = 12'h000;
rom[418] = 12'h00f;
rom[419] = 12'h00f;
rom[420] = 12'h00f;
rom[421] = 12'h00f;
rom[422] = 12'h00f;
rom[423] = 12'h00f;
rom[424] = 12'h000;
rom[425] = 12'h000;
rom[426] = 12'h000;
rom[427] = 12'h000;
rom[428] = 12'h000;
rom[429] = 12'h000;
rom[430] = 12'h000;
rom[431] = 12'h000;
rom[432] = 12'h000;
rom[433] = 12'h000;
rom[434] = 12'h00f;
rom[435] = 12'h00f;
rom[436] = 12'h00f;
rom[437] = 12'h00f;
rom[438] = 12'h00f;
rom[439] = 12'h00f;
rom[440] = 12'h000;
rom[441] = 12'h000;
rom[442] = 12'h000;
rom[443] = 12'h000;
rom[444] = 12'h00f;
rom[445] = 12'h00f;
rom[446] = 12'h00f;
rom[447] = 12'h00f;
rom[448] = 12'h00f;
rom[449] = 12'h00f;
rom[450] = 12'h000;
rom[451] = 12'h000;
rom[452] = 12'h000;
rom[453] = 12'h000;
rom[454] = 12'h000;
rom[455] = 12'h000;
rom[456] = 12'h000;
rom[457] = 12'h000;
rom[458] = 12'h000;
rom[459] = 12'h000;
rom[460] = 12'h00f;
rom[461] = 12'h00f;
rom[462] = 12'h00f;
rom[463] = 12'h00f;
rom[464] = 12'h00f;
rom[465] = 12'h00f;
rom[466] = 12'h000;
rom[467] = 12'h000;
rom[468] = 12'h000;
rom[469] = 12'h000;
rom[470] = 12'h00f;
rom[471] = 12'h00f;
rom[472] = 12'h00f;
rom[473] = 12'h00f;
rom[474] = 12'h000;
rom[475] = 12'h000;
rom[476] = 12'h000;
rom[477] = 12'h000;
rom[478] = 12'h000;
rom[479] = 12'h000;
rom[480] = 12'h000;
rom[481] = 12'h000;
rom[482] = 12'h000;
rom[483] = 12'h000;
rom[484] = 12'h000;
rom[485] = 12'h000;
rom[486] = 12'h000;
rom[487] = 12'h000;
rom[488] = 12'h00f;
rom[489] = 12'h00f;
rom[490] = 12'h00f;
rom[491] = 12'h00f;
rom[492] = 12'h000;
rom[493] = 12'h000;
rom[494] = 12'h000;
rom[495] = 12'h000;
rom[496] = 12'h00f;
rom[497] = 12'h00f;
rom[498] = 12'h00f;
rom[499] = 12'h00f;
rom[500] = 12'h000;
rom[501] = 12'h000;
rom[502] = 12'h000;
rom[503] = 12'h000;
rom[504] = 12'h000;
rom[505] = 12'h000;
rom[506] = 12'h000;
rom[507] = 12'h000;
rom[508] = 12'h000;
rom[509] = 12'h000;
rom[510] = 12'h000;
rom[511] = 12'h000;
rom[512] = 12'h000;
rom[513] = 12'h000;
rom[514] = 12'h00f;
rom[515] = 12'h00f;
rom[516] = 12'h00f;
rom[517] = 12'h00f;
rom[518] = 12'h000;
rom[519] = 12'h000;
rom[520] = 12'h000;
rom[521] = 12'h000;
rom[522] = 12'h00f;
rom[523] = 12'h00f;
rom[524] = 12'h000;
rom[525] = 12'h000;
rom[526] = 12'h000;
rom[527] = 12'h000;
rom[528] = 12'h007;
rom[529] = 12'h007;
rom[530] = 12'h000;
rom[531] = 12'h000;
rom[532] = 12'h007;
rom[533] = 12'h007;
rom[534] = 12'h000;
rom[535] = 12'h000;
rom[536] = 12'h007;
rom[537] = 12'h007;
rom[538] = 12'h000;
rom[539] = 12'h000;
rom[540] = 12'h000;
rom[541] = 12'h000;
rom[542] = 12'h00f;
rom[543] = 12'h00f;
rom[544] = 12'h000;
rom[545] = 12'h000;
rom[546] = 12'h000;
rom[547] = 12'h000;
rom[548] = 12'h00f;
rom[549] = 12'h00f;
rom[550] = 12'h000;
rom[551] = 12'h000;
rom[552] = 12'h000;
rom[553] = 12'h000;
rom[554] = 12'h007;
rom[555] = 12'h007;
rom[556] = 12'h000;
rom[557] = 12'h000;
rom[558] = 12'h007;
rom[559] = 12'h007;
rom[560] = 12'h000;
rom[561] = 12'h000;
rom[562] = 12'h007;
rom[563] = 12'h007;
rom[564] = 12'h000;
rom[565] = 12'h000;
rom[566] = 12'h000;
rom[567] = 12'h000;
rom[568] = 12'h00f;
rom[569] = 12'h00f;
rom[570] = 12'h000;
rom[571] = 12'h000;
rom[572] = 12'h000;
rom[573] = 12'h000;
rom[574] = 12'h000;
rom[575] = 12'h000;
rom[576] = 12'h000;
rom[577] = 12'h000;
rom[578] = 12'h007;
rom[579] = 12'h007;
rom[580] = 12'h000;
rom[581] = 12'h000;
rom[582] = 12'h007;
rom[583] = 12'h007;
rom[584] = 12'h000;
rom[585] = 12'h000;
rom[586] = 12'h007;
rom[587] = 12'h007;
rom[588] = 12'h000;
rom[589] = 12'h000;
rom[590] = 12'h007;
rom[591] = 12'h007;
rom[592] = 12'h000;
rom[593] = 12'h000;
rom[594] = 12'h000;
rom[595] = 12'h000;
rom[596] = 12'h000;
rom[597] = 12'h000;
rom[598] = 12'h000;
rom[599] = 12'h000;
rom[600] = 12'h000;
rom[601] = 12'h000;
rom[602] = 12'h000;
rom[603] = 12'h000;
rom[604] = 12'h007;
rom[605] = 12'h007;
rom[606] = 12'h000;
rom[607] = 12'h000;
rom[608] = 12'h007;
rom[609] = 12'h007;
rom[610] = 12'h000;
rom[611] = 12'h000;
rom[612] = 12'h007;
rom[613] = 12'h007;
rom[614] = 12'h000;
rom[615] = 12'h000;
rom[616] = 12'h007;
rom[617] = 12'h007;
rom[618] = 12'h000;
rom[619] = 12'h000;
rom[620] = 12'h000;
rom[621] = 12'h000;
rom[622] = 12'h000;
rom[623] = 12'h000;
rom[624] = 12'h000;
rom[625] = 12'h000;
rom[626] = 12'h00f;
rom[627] = 12'h00f;
rom[628] = 12'h000;
rom[629] = 12'h000;
rom[630] = 12'h000;
rom[631] = 12'h000;
rom[632] = 12'h007;
rom[633] = 12'h007;
rom[634] = 12'h000;
rom[635] = 12'h000;
rom[636] = 12'h007;
rom[637] = 12'h007;
rom[638] = 12'h000;
rom[639] = 12'h000;
rom[640] = 12'h007;
rom[641] = 12'h007;
rom[642] = 12'h000;
rom[643] = 12'h000;
rom[644] = 12'h000;
rom[645] = 12'h000;
rom[646] = 12'h00f;
rom[647] = 12'h00f;
rom[648] = 12'h000;
rom[649] = 12'h000;
rom[650] = 12'h000;
rom[651] = 12'h000;
rom[652] = 12'h00f;
rom[653] = 12'h00f;
rom[654] = 12'h000;
rom[655] = 12'h000;
rom[656] = 12'h000;
rom[657] = 12'h000;
rom[658] = 12'h007;
rom[659] = 12'h007;
rom[660] = 12'h000;
rom[661] = 12'h000;
rom[662] = 12'h007;
rom[663] = 12'h007;
rom[664] = 12'h000;
rom[665] = 12'h000;
rom[666] = 12'h007;
rom[667] = 12'h007;
rom[668] = 12'h000;
rom[669] = 12'h000;
rom[670] = 12'h000;
rom[671] = 12'h000;
rom[672] = 12'h00f;
rom[673] = 12'h00f;
rom[674] = 12'h000;
rom[675] = 12'h000;
rom[676] = 12'h000;
rom[677] = 12'h000;
rom[678] = 12'h00f;
rom[679] = 12'h00f;
rom[680] = 12'h00f;
rom[681] = 12'h00f;
rom[682] = 12'h000;
rom[683] = 12'h000;
rom[684] = 12'h000;
rom[685] = 12'h000;
rom[686] = 12'h000;
rom[687] = 12'h000;
rom[688] = 12'h000;
rom[689] = 12'h000;
rom[690] = 12'h000;
rom[691] = 12'h000;
rom[692] = 12'h000;
rom[693] = 12'h000;
rom[694] = 12'h000;
rom[695] = 12'h000;
rom[696] = 12'h00f;
rom[697] = 12'h00f;
rom[698] = 12'h00f;
rom[699] = 12'h00f;
rom[700] = 12'h000;
rom[701] = 12'h000;
rom[702] = 12'h000;
rom[703] = 12'h000;
rom[704] = 12'h00f;
rom[705] = 12'h00f;
rom[706] = 12'h00f;
rom[707] = 12'h00f;
rom[708] = 12'h000;
rom[709] = 12'h000;
rom[710] = 12'h000;
rom[711] = 12'h000;
rom[712] = 12'h000;
rom[713] = 12'h000;
rom[714] = 12'h000;
rom[715] = 12'h000;
rom[716] = 12'h000;
rom[717] = 12'h000;
rom[718] = 12'h000;
rom[719] = 12'h000;
rom[720] = 12'h000;
rom[721] = 12'h000;
rom[722] = 12'h00f;
rom[723] = 12'h00f;
rom[724] = 12'h00f;
rom[725] = 12'h00f;
rom[726] = 12'h000;
rom[727] = 12'h000;
rom[728] = 12'h000;
rom[729] = 12'h000;
rom[730] = 12'h00f;
rom[731] = 12'h00f;
rom[732] = 12'h00f;
rom[733] = 12'h00f;
rom[734] = 12'h00f;
rom[735] = 12'h00f;
rom[736] = 12'h000;
rom[737] = 12'h000;
rom[738] = 12'h000;
rom[739] = 12'h000;
rom[740] = 12'h000;
rom[741] = 12'h000;
rom[742] = 12'h000;
rom[743] = 12'h000;
rom[744] = 12'h000;
rom[745] = 12'h000;
rom[746] = 12'h00f;
rom[747] = 12'h00f;
rom[748] = 12'h00f;
rom[749] = 12'h00f;
rom[750] = 12'h00f;
rom[751] = 12'h00f;
rom[752] = 12'h000;
rom[753] = 12'h000;
rom[754] = 12'h000;
rom[755] = 12'h000;
rom[756] = 12'h00f;
rom[757] = 12'h00f;
rom[758] = 12'h00f;
rom[759] = 12'h00f;
rom[760] = 12'h00f;
rom[761] = 12'h00f;
rom[762] = 12'h000;
rom[763] = 12'h000;
rom[764] = 12'h000;
rom[765] = 12'h000;
rom[766] = 12'h000;
rom[767] = 12'h000;
rom[768] = 12'h000;
rom[769] = 12'h000;
rom[770] = 12'h000;
rom[771] = 12'h000;
rom[772] = 12'h00f;
rom[773] = 12'h00f;
rom[774] = 12'h00f;
rom[775] = 12'h00f;
rom[776] = 12'h00f;
rom[777] = 12'h00f;
rom[778] = 12'h000;
rom[779] = 12'h000;
rom[780] = 12'h000;
rom[781] = 12'h000;
rom[782] = 12'h00f;
rom[783] = 12'h00f;
rom[784] = 12'h00f;
rom[785] = 12'h00f;
rom[786] = 12'h00f;
rom[787] = 12'h00f;
rom[788] = 12'h000;
rom[789] = 12'h000;
rom[790] = 12'h000;
rom[791] = 12'h000;
rom[792] = 12'h000;
rom[793] = 12'h000;
rom[794] = 12'h000;
rom[795] = 12'h000;
rom[796] = 12'h000;
rom[797] = 12'h000;
rom[798] = 12'h00f;
rom[799] = 12'h00f;
rom[800] = 12'h00f;
rom[801] = 12'h00f;
rom[802] = 12'h00f;
rom[803] = 12'h00f;
rom[804] = 12'h000;
rom[805] = 12'h000;
rom[806] = 12'h000;
rom[807] = 12'h000;
rom[808] = 12'h00f;
rom[809] = 12'h00f;
rom[810] = 12'h00f;
rom[811] = 12'h00f;
rom[812] = 12'h00f;
rom[813] = 12'h00f;
rom[814] = 12'h000;
rom[815] = 12'h000;
rom[816] = 12'h000;
rom[817] = 12'h000;
rom[818] = 12'h000;
rom[819] = 12'h000;
rom[820] = 12'h000;
rom[821] = 12'h000;
rom[822] = 12'h000;
rom[823] = 12'h000;
rom[824] = 12'h00f;
rom[825] = 12'h00f;
rom[826] = 12'h00f;
rom[827] = 12'h00f;
rom[828] = 12'h00f;
rom[829] = 12'h00f;
rom[830] = 12'h000;
rom[831] = 12'h000;
rom[832] = 12'h000;
rom[833] = 12'h000;
rom[834] = 12'h00f;
rom[835] = 12'h00f;
rom[836] = 12'h00f;
rom[837] = 12'h00f;
rom[838] = 12'h00f;
rom[839] = 12'h00f;
rom[840] = 12'h000;
rom[841] = 12'h000;
rom[842] = 12'h000;
rom[843] = 12'h000;
rom[844] = 12'h000;
rom[845] = 12'h000;
rom[846] = 12'h000;
rom[847] = 12'h000;
rom[848] = 12'h000;
rom[849] = 12'h000;
rom[850] = 12'h00f;
rom[851] = 12'h00f;
rom[852] = 12'h00f;
rom[853] = 12'h00f;
rom[854] = 12'h00f;
rom[855] = 12'h00f;
rom[856] = 12'h000;
rom[857] = 12'h000;
rom[858] = 12'h000;
rom[859] = 12'h000;
rom[860] = 12'h00f;
rom[861] = 12'h00f;
rom[862] = 12'h00f;
rom[863] = 12'h00f;
rom[864] = 12'h00f;
rom[865] = 12'h00f;
rom[866] = 12'h000;
rom[867] = 12'h000;
rom[868] = 12'h000;
rom[869] = 12'h000;
rom[870] = 12'h000;
rom[871] = 12'h000;
rom[872] = 12'h000;
rom[873] = 12'h000;
rom[874] = 12'h000;
rom[875] = 12'h000;
rom[876] = 12'h00f;
rom[877] = 12'h00f;
rom[878] = 12'h00f;
rom[879] = 12'h00f;
rom[880] = 12'h00f;
rom[881] = 12'h00f;
rom[882] = 12'h000;
rom[883] = 12'h000;
rom[884] = 12'h000;
rom[885] = 12'h000;
rom[886] = 12'h00f;
rom[887] = 12'h00f;
rom[888] = 12'h00f;
rom[889] = 12'h00f;
rom[890] = 12'h00f;
rom[891] = 12'h00f;
rom[892] = 12'h000;
rom[893] = 12'h000;
rom[894] = 12'h000;
rom[895] = 12'h000;
rom[896] = 12'h000;
rom[897] = 12'h000;
rom[898] = 12'h000;
rom[899] = 12'h000;
rom[900] = 12'h000;
rom[901] = 12'h000;
rom[902] = 12'h00f;
rom[903] = 12'h00f;
rom[904] = 12'h00f;
rom[905] = 12'h00f;
rom[906] = 12'h00f;
rom[907] = 12'h00f;
rom[908] = 12'h000;
rom[909] = 12'h000;
rom[910] = 12'h000;
rom[911] = 12'h000;
rom[912] = 12'h00f;
rom[913] = 12'h00f;
rom[914] = 12'h00f;
rom[915] = 12'h00f;
rom[916] = 12'h00f;
rom[917] = 12'h00f;
rom[918] = 12'h000;
rom[919] = 12'h000;
rom[920] = 12'h000;
rom[921] = 12'h000;
rom[922] = 12'h000;
rom[923] = 12'h000;
rom[924] = 12'h000;
rom[925] = 12'h000;
rom[926] = 12'h000;
rom[927] = 12'h000;
rom[928] = 12'h00f;
rom[929] = 12'h00f;
rom[930] = 12'h00f;
rom[931] = 12'h00f;
rom[932] = 12'h00f;
rom[933] = 12'h00f;
rom[934] = 12'h000;
rom[935] = 12'h000;
rom[936] = 12'h000;
rom[937] = 12'h000;
rom[938] = 12'h00f;
rom[939] = 12'h00f;
rom[940] = 12'h00f;
rom[941] = 12'h00f;
rom[942] = 12'h00f;
rom[943] = 12'h00f;
rom[944] = 12'h000;
rom[945] = 12'h000;
rom[946] = 12'h000;
rom[947] = 12'h000;
rom[948] = 12'h000;
rom[949] = 12'h000;
rom[950] = 12'h000;
rom[951] = 12'h000;
rom[952] = 12'h000;
rom[953] = 12'h000;
rom[954] = 12'h00f;
rom[955] = 12'h00f;
rom[956] = 12'h00f;
rom[957] = 12'h00f;
rom[958] = 12'h00f;
rom[959] = 12'h00f;
rom[960] = 12'h000;
rom[961] = 12'h000;
rom[962] = 12'h000;
rom[963] = 12'h000;
rom[964] = 12'h00f;
rom[965] = 12'h00f;
rom[966] = 12'h00f;
rom[967] = 12'h00f;
rom[968] = 12'h00f;
rom[969] = 12'h00f;
rom[970] = 12'h000;
rom[971] = 12'h000;
rom[972] = 12'h000;
rom[973] = 12'h000;
rom[974] = 12'h000;
rom[975] = 12'h000;
rom[976] = 12'h000;
rom[977] = 12'h000;
rom[978] = 12'h000;
rom[979] = 12'h000;
rom[980] = 12'h00f;
rom[981] = 12'h00f;
rom[982] = 12'h00f;
rom[983] = 12'h00f;
rom[984] = 12'h00f;
rom[985] = 12'h00f;
rom[986] = 12'h000;
rom[987] = 12'h000;
rom[988] = 12'h000;
rom[989] = 12'h000;
rom[990] = 12'h00f;
rom[991] = 12'h00f;
rom[992] = 12'h00f;
rom[993] = 12'h00f;
rom[994] = 12'h000;
rom[995] = 12'h000;
rom[996] = 12'h00f;
rom[997] = 12'h00f;
rom[998] = 12'h00f;
rom[999] = 12'h00f;
rom[1000] = 12'h00f;
rom[1001] = 12'h00f;
rom[1002] = 12'h00f;
rom[1003] = 12'h00f;
rom[1004] = 12'h00f;
rom[1005] = 12'h00f;
rom[1006] = 12'h000;
rom[1007] = 12'h000;
rom[1008] = 12'h00f;
rom[1009] = 12'h00f;
rom[1010] = 12'h00f;
rom[1011] = 12'h00f;
rom[1012] = 12'h000;
rom[1013] = 12'h000;
rom[1014] = 12'h000;
rom[1015] = 12'h000;
rom[1016] = 12'h00f;
rom[1017] = 12'h00f;
rom[1018] = 12'h00f;
rom[1019] = 12'h00f;
rom[1020] = 12'h000;
rom[1021] = 12'h000;
rom[1022] = 12'h00f;
rom[1023] = 12'h00f;
rom[1024] = 12'h00f;
rom[1025] = 12'h00f;
rom[1026] = 12'h00f;
rom[1027] = 12'h00f;
rom[1028] = 12'h00f;
rom[1029] = 12'h00f;
rom[1030] = 12'h00f;
rom[1031] = 12'h00f;
rom[1032] = 12'h000;
rom[1033] = 12'h000;
rom[1034] = 12'h00f;
rom[1035] = 12'h00f;
rom[1036] = 12'h00f;
rom[1037] = 12'h00f;
rom[1038] = 12'h000;
rom[1039] = 12'h000;
rom[1040] = 12'h000;
rom[1041] = 12'h000;
rom[1042] = 12'h00f;
rom[1043] = 12'h00f;
rom[1044] = 12'h000;
rom[1045] = 12'h000;
rom[1046] = 12'h00f;
rom[1047] = 12'h00f;
rom[1048] = 12'h00f;
rom[1049] = 12'h00f;
rom[1050] = 12'h00f;
rom[1051] = 12'h00f;
rom[1052] = 12'h00f;
rom[1053] = 12'h00f;
rom[1054] = 12'h00f;
rom[1055] = 12'h00f;
rom[1056] = 12'h00f;
rom[1057] = 12'h00f;
rom[1058] = 12'h00f;
rom[1059] = 12'h00f;
rom[1060] = 12'h000;
rom[1061] = 12'h000;
rom[1062] = 12'h00f;
rom[1063] = 12'h00f;
rom[1064] = 12'h000;
rom[1065] = 12'h000;
rom[1066] = 12'h000;
rom[1067] = 12'h000;
rom[1068] = 12'h00f;
rom[1069] = 12'h00f;
rom[1070] = 12'h000;
rom[1071] = 12'h000;
rom[1072] = 12'h00f;
rom[1073] = 12'h00f;
rom[1074] = 12'h00f;
rom[1075] = 12'h00f;
rom[1076] = 12'h00f;
rom[1077] = 12'h00f;
rom[1078] = 12'h00f;
rom[1079] = 12'h00f;
rom[1080] = 12'h00f;
rom[1081] = 12'h00f;
rom[1082] = 12'h00f;
rom[1083] = 12'h00f;
rom[1084] = 12'h00f;
rom[1085] = 12'h00f;
rom[1086] = 12'h000;
rom[1087] = 12'h000;
rom[1088] = 12'h00f;
rom[1089] = 12'h00f;
rom[1090] = 12'h000;
rom[1091] = 12'h000;
rom[1092] = 12'h000;
rom[1093] = 12'h000;
rom[1094] = 12'h000;
rom[1095] = 12'h000;
rom[1096] = 12'h00f;
rom[1097] = 12'h00f;
rom[1098] = 12'h00f;
rom[1099] = 12'h00f;
rom[1100] = 12'h00f;
rom[1101] = 12'h00f;
rom[1102] = 12'h00f;
rom[1103] = 12'h00f;
rom[1104] = 12'h00f;
rom[1105] = 12'h00f;
rom[1106] = 12'h00f;
rom[1107] = 12'h00f;
rom[1108] = 12'h00f;
rom[1109] = 12'h00f;
rom[1110] = 12'h00f;
rom[1111] = 12'h00f;
rom[1112] = 12'h00f;
rom[1113] = 12'h00f;
rom[1114] = 12'h000;
rom[1115] = 12'h000;
rom[1116] = 12'h000;
rom[1117] = 12'h000;
rom[1118] = 12'h000;
rom[1119] = 12'h000;
rom[1120] = 12'h000;
rom[1121] = 12'h000;
rom[1122] = 12'h00f;
rom[1123] = 12'h00f;
rom[1124] = 12'h00f;
rom[1125] = 12'h00f;
rom[1126] = 12'h00f;
rom[1127] = 12'h00f;
rom[1128] = 12'h00f;
rom[1129] = 12'h00f;
rom[1130] = 12'h00f;
rom[1131] = 12'h00f;
rom[1132] = 12'h00f;
rom[1133] = 12'h00f;
rom[1134] = 12'h00f;
rom[1135] = 12'h00f;
rom[1136] = 12'h00f;
rom[1137] = 12'h00f;
rom[1138] = 12'h00f;
rom[1139] = 12'h00f;
rom[1140] = 12'h000;
rom[1141] = 12'h000;
rom[1142] = 12'h000;
rom[1143] = 12'h000;
rom[1144] = 12'h000;
rom[1145] = 12'h000;
rom[1146] = 12'h000;
rom[1147] = 12'h000;
rom[1148] = 12'h000;
rom[1149] = 12'h000;
rom[1150] = 12'h000;
rom[1151] = 12'h000;
rom[1152] = 12'h000;
rom[1153] = 12'h000;
rom[1154] = 12'h000;
rom[1155] = 12'h000;
rom[1156] = 12'h000;
rom[1157] = 12'h000;
rom[1158] = 12'h000;
rom[1159] = 12'h000;
rom[1160] = 12'h000;
rom[1161] = 12'h000;
rom[1162] = 12'h000;
rom[1163] = 12'h000;
rom[1164] = 12'h000;
rom[1165] = 12'h000;
rom[1166] = 12'h000;
rom[1167] = 12'h000;
rom[1168] = 12'h000;
rom[1169] = 12'h000;
rom[1170] = 12'h000;
rom[1171] = 12'h000;
rom[1172] = 12'h000;
rom[1173] = 12'h000;
rom[1174] = 12'h000;
rom[1175] = 12'h000;
rom[1176] = 12'h000;
rom[1177] = 12'h000;
rom[1178] = 12'h000;
rom[1179] = 12'h000;
rom[1180] = 12'h000;
rom[1181] = 12'h000;
rom[1182] = 12'h000;
rom[1183] = 12'h000;
rom[1184] = 12'h000;
rom[1185] = 12'h000;
rom[1186] = 12'h000;
rom[1187] = 12'h000;
rom[1188] = 12'h000;
rom[1189] = 12'h000;
rom[1190] = 12'h000;
rom[1191] = 12'h000;
rom[1192] = 12'h000;
rom[1193] = 12'h000;
rom[1194] = 12'h000;
rom[1195] = 12'h000;
  end
  endmodule

    module one_rom (                       //один
  input  wire    [13:0]     addr,
  output wire    [11:0]     word
);

  logic [11:0] rom [(46 * 26)];

  assign word = rom[addr];

  initial begin
rom[0] = 12'h000;
rom[1] = 12'h000;
rom[2] = 12'h000;
rom[3] = 12'h000;
rom[4] = 12'h000;
rom[5] = 12'h000;
rom[6] = 12'h000;
rom[7] = 12'h000;
rom[8] = 12'h000;
rom[9] = 12'h000;
rom[10] = 12'h000;
rom[11] = 12'h000;
rom[12] = 12'h000;
rom[13] = 12'h000;
rom[14] = 12'h000;
rom[15] = 12'h000;
rom[16] = 12'h000;
rom[17] = 12'h000;
rom[18] = 12'h000;
rom[19] = 12'h000;
rom[20] = 12'h000;
rom[21] = 12'h000;
rom[22] = 12'h000;
rom[23] = 12'h000;
rom[24] = 12'h000;
rom[25] = 12'h000;
rom[26] = 12'h000;
rom[27] = 12'h000;
rom[28] = 12'h000;
rom[29] = 12'h000;
rom[30] = 12'h000;
rom[31] = 12'h000;
rom[32] = 12'h000;
rom[33] = 12'h000;
rom[34] = 12'h000;
rom[35] = 12'h000;
rom[36] = 12'h000;
rom[37] = 12'h000;
rom[38] = 12'h000;
rom[39] = 12'h000;
rom[40] = 12'h000;
rom[41] = 12'h000;
rom[42] = 12'h000;
rom[43] = 12'h000;
rom[44] = 12'h000;
rom[45] = 12'h000;
rom[46] = 12'h000;
rom[47] = 12'h000;
rom[48] = 12'h000;
rom[49] = 12'h000;
rom[50] = 12'h000;
rom[51] = 12'h000;
rom[52] = 12'h000;
rom[53] = 12'h000;
rom[54] = 12'h000;
rom[55] = 12'h000;
rom[56] = 12'h000;
rom[57] = 12'h000;
rom[58] = 12'h007;
rom[59] = 12'h007;
rom[60] = 12'h000;
rom[61] = 12'h000;
rom[62] = 12'h007;
rom[63] = 12'h007;
rom[64] = 12'h000;
rom[65] = 12'h000;
rom[66] = 12'h007;
rom[67] = 12'h007;
rom[68] = 12'h000;
rom[69] = 12'h000;
rom[70] = 12'h007;
rom[71] = 12'h007;
rom[72] = 12'h000;
rom[73] = 12'h000;
rom[74] = 12'h000;
rom[75] = 12'h000;
rom[76] = 12'h000;
rom[77] = 12'h000;
rom[78] = 12'h000;
rom[79] = 12'h000;
rom[80] = 12'h000;
rom[81] = 12'h000;
rom[82] = 12'h000;
rom[83] = 12'h000;
rom[84] = 12'h007;
rom[85] = 12'h007;
rom[86] = 12'h000;
rom[87] = 12'h000;
rom[88] = 12'h007;
rom[89] = 12'h007;
rom[90] = 12'h000;
rom[91] = 12'h000;
rom[92] = 12'h007;
rom[93] = 12'h007;
rom[94] = 12'h000;
rom[95] = 12'h000;
rom[96] = 12'h007;
rom[97] = 12'h007;
rom[98] = 12'h000;
rom[99] = 12'h000;
rom[100] = 12'h000;
rom[101] = 12'h000;
rom[102] = 12'h000;
rom[103] = 12'h000;
rom[104] = 12'h000;
rom[105] = 12'h000;
rom[106] = 12'h007;
rom[107] = 12'h007;
rom[108] = 12'h000;
rom[109] = 12'h000;
rom[110] = 12'h000;
rom[111] = 12'h000;
rom[112] = 12'h007;
rom[113] = 12'h007;
rom[114] = 12'h000;
rom[115] = 12'h000;
rom[116] = 12'h007;
rom[117] = 12'h007;
rom[118] = 12'h000;
rom[119] = 12'h000;
rom[120] = 12'h007;
rom[121] = 12'h007;
rom[122] = 12'h000;
rom[123] = 12'h000;
rom[124] = 12'h000;
rom[125] = 12'h000;
rom[126] = 12'h00f;
rom[127] = 12'h00f;
rom[128] = 12'h000;
rom[129] = 12'h000;
rom[130] = 12'h000;
rom[131] = 12'h000;
rom[132] = 12'h007;
rom[133] = 12'h007;
rom[134] = 12'h000;
rom[135] = 12'h000;
rom[136] = 12'h000;
rom[137] = 12'h000;
rom[138] = 12'h007;
rom[139] = 12'h007;
rom[140] = 12'h000;
rom[141] = 12'h000;
rom[142] = 12'h007;
rom[143] = 12'h007;
rom[144] = 12'h000;
rom[145] = 12'h000;
rom[146] = 12'h007;
rom[147] = 12'h007;
rom[148] = 12'h000;
rom[149] = 12'h000;
rom[150] = 12'h000;
rom[151] = 12'h000;
rom[152] = 12'h00f;
rom[153] = 12'h00f;
rom[154] = 12'h000;
rom[155] = 12'h000;
rom[156] = 12'h000;
rom[157] = 12'h000;
rom[158] = 12'h000;
rom[159] = 12'h000;
rom[160] = 12'h007;
rom[161] = 12'h007;
rom[162] = 12'h000;
rom[163] = 12'h000;
rom[164] = 12'h000;
rom[165] = 12'h000;
rom[166] = 12'h007;
rom[167] = 12'h007;
rom[168] = 12'h000;
rom[169] = 12'h000;
rom[170] = 12'h007;
rom[171] = 12'h007;
rom[172] = 12'h000;
rom[173] = 12'h000;
rom[174] = 12'h000;
rom[175] = 12'h000;
rom[176] = 12'h00f;
rom[177] = 12'h00f;
rom[178] = 12'h00f;
rom[179] = 12'h00f;
rom[180] = 12'h000;
rom[181] = 12'h000;
rom[182] = 12'h000;
rom[183] = 12'h000;
rom[184] = 12'h000;
rom[185] = 12'h000;
rom[186] = 12'h007;
rom[187] = 12'h007;
rom[188] = 12'h000;
rom[189] = 12'h000;
rom[190] = 12'h000;
rom[191] = 12'h000;
rom[192] = 12'h007;
rom[193] = 12'h007;
rom[194] = 12'h000;
rom[195] = 12'h000;
rom[196] = 12'h007;
rom[197] = 12'h007;
rom[198] = 12'h000;
rom[199] = 12'h000;
rom[200] = 12'h000;
rom[201] = 12'h000;
rom[202] = 12'h00f;
rom[203] = 12'h00f;
rom[204] = 12'h00f;
rom[205] = 12'h00f;
rom[206] = 12'h000;
rom[207] = 12'h000;
rom[208] = 12'h000;
rom[209] = 12'h000;
rom[210] = 12'h007;
rom[211] = 12'h007;
rom[212] = 12'h000;
rom[213] = 12'h000;
rom[214] = 12'h007;
rom[215] = 12'h007;
rom[216] = 12'h000;
rom[217] = 12'h000;
rom[218] = 12'h000;
rom[219] = 12'h000;
rom[220] = 12'h000;
rom[221] = 12'h000;
rom[222] = 12'h000;
rom[223] = 12'h000;
rom[224] = 12'h000;
rom[225] = 12'h000;
rom[226] = 12'h00f;
rom[227] = 12'h00f;
rom[228] = 12'h00f;
rom[229] = 12'h00f;
rom[230] = 12'h00f;
rom[231] = 12'h00f;
rom[232] = 12'h000;
rom[233] = 12'h000;
rom[234] = 12'h000;
rom[235] = 12'h000;
rom[236] = 12'h007;
rom[237] = 12'h007;
rom[238] = 12'h000;
rom[239] = 12'h000;
rom[240] = 12'h007;
rom[241] = 12'h007;
rom[242] = 12'h000;
rom[243] = 12'h000;
rom[244] = 12'h000;
rom[245] = 12'h000;
rom[246] = 12'h000;
rom[247] = 12'h000;
rom[248] = 12'h000;
rom[249] = 12'h000;
rom[250] = 12'h000;
rom[251] = 12'h000;
rom[252] = 12'h00f;
rom[253] = 12'h00f;
rom[254] = 12'h00f;
rom[255] = 12'h00f;
rom[256] = 12'h00f;
rom[257] = 12'h00f;
rom[258] = 12'h000;
rom[259] = 12'h000;
rom[260] = 12'h000;
rom[261] = 12'h000;
rom[262] = 12'h000;
rom[263] = 12'h000;
rom[264] = 12'h007;
rom[265] = 12'h007;
rom[266] = 12'h000;
rom[267] = 12'h000;
rom[268] = 12'h000;
rom[269] = 12'h000;
rom[270] = 12'h000;
rom[271] = 12'h000;
rom[272] = 12'h000;
rom[273] = 12'h000;
rom[274] = 12'h000;
rom[275] = 12'h000;
rom[276] = 12'h000;
rom[277] = 12'h000;
rom[278] = 12'h00f;
rom[279] = 12'h00f;
rom[280] = 12'h00f;
rom[281] = 12'h00f;
rom[282] = 12'h00f;
rom[283] = 12'h00f;
rom[284] = 12'h000;
rom[285] = 12'h000;
rom[286] = 12'h000;
rom[287] = 12'h000;
rom[288] = 12'h000;
rom[289] = 12'h000;
rom[290] = 12'h007;
rom[291] = 12'h007;
rom[292] = 12'h000;
rom[293] = 12'h000;
rom[294] = 12'h000;
rom[295] = 12'h000;
rom[296] = 12'h000;
rom[297] = 12'h000;
rom[298] = 12'h000;
rom[299] = 12'h000;
rom[300] = 12'h000;
rom[301] = 12'h000;
rom[302] = 12'h000;
rom[303] = 12'h000;
rom[304] = 12'h00f;
rom[305] = 12'h00f;
rom[306] = 12'h00f;
rom[307] = 12'h00f;
rom[308] = 12'h00f;
rom[309] = 12'h00f;
rom[310] = 12'h000;
rom[311] = 12'h000;
rom[312] = 12'h000;
rom[313] = 12'h000;
rom[314] = 12'h007;
rom[315] = 12'h007;
rom[316] = 12'h000;
rom[317] = 12'h000;
rom[318] = 12'h007;
rom[319] = 12'h007;
rom[320] = 12'h000;
rom[321] = 12'h000;
rom[322] = 12'h000;
rom[323] = 12'h000;
rom[324] = 12'h000;
rom[325] = 12'h000;
rom[326] = 12'h000;
rom[327] = 12'h000;
rom[328] = 12'h000;
rom[329] = 12'h000;
rom[330] = 12'h00f;
rom[331] = 12'h00f;
rom[332] = 12'h00f;
rom[333] = 12'h00f;
rom[334] = 12'h00f;
rom[335] = 12'h00f;
rom[336] = 12'h000;
rom[337] = 12'h000;
rom[338] = 12'h000;
rom[339] = 12'h000;
rom[340] = 12'h007;
rom[341] = 12'h007;
rom[342] = 12'h000;
rom[343] = 12'h000;
rom[344] = 12'h007;
rom[345] = 12'h007;
rom[346] = 12'h000;
rom[347] = 12'h000;
rom[348] = 12'h000;
rom[349] = 12'h000;
rom[350] = 12'h000;
rom[351] = 12'h000;
rom[352] = 12'h000;
rom[353] = 12'h000;
rom[354] = 12'h000;
rom[355] = 12'h000;
rom[356] = 12'h00f;
rom[357] = 12'h00f;
rom[358] = 12'h00f;
rom[359] = 12'h00f;
rom[360] = 12'h00f;
rom[361] = 12'h00f;
rom[362] = 12'h000;
rom[363] = 12'h000;
rom[364] = 12'h000;
rom[365] = 12'h000;
rom[366] = 12'h000;
rom[367] = 12'h000;
rom[368] = 12'h007;
rom[369] = 12'h007;
rom[370] = 12'h000;
rom[371] = 12'h000;
rom[372] = 12'h000;
rom[373] = 12'h000;
rom[374] = 12'h000;
rom[375] = 12'h000;
rom[376] = 12'h000;
rom[377] = 12'h000;
rom[378] = 12'h000;
rom[379] = 12'h000;
rom[380] = 12'h000;
rom[381] = 12'h000;
rom[382] = 12'h00f;
rom[383] = 12'h00f;
rom[384] = 12'h00f;
rom[385] = 12'h00f;
rom[386] = 12'h00f;
rom[387] = 12'h00f;
rom[388] = 12'h000;
rom[389] = 12'h000;
rom[390] = 12'h000;
rom[391] = 12'h000;
rom[392] = 12'h000;
rom[393] = 12'h000;
rom[394] = 12'h007;
rom[395] = 12'h007;
rom[396] = 12'h000;
rom[397] = 12'h000;
rom[398] = 12'h000;
rom[399] = 12'h000;
rom[400] = 12'h000;
rom[401] = 12'h000;
rom[402] = 12'h000;
rom[403] = 12'h000;
rom[404] = 12'h000;
rom[405] = 12'h000;
rom[406] = 12'h000;
rom[407] = 12'h000;
rom[408] = 12'h00f;
rom[409] = 12'h00f;
rom[410] = 12'h00f;
rom[411] = 12'h00f;
rom[412] = 12'h00f;
rom[413] = 12'h00f;
rom[414] = 12'h000;
rom[415] = 12'h000;
rom[416] = 12'h000;
rom[417] = 12'h000;
rom[418] = 12'h007;
rom[419] = 12'h007;
rom[420] = 12'h000;
rom[421] = 12'h000;
rom[422] = 12'h007;
rom[423] = 12'h007;
rom[424] = 12'h000;
rom[425] = 12'h000;
rom[426] = 12'h000;
rom[427] = 12'h000;
rom[428] = 12'h000;
rom[429] = 12'h000;
rom[430] = 12'h000;
rom[431] = 12'h000;
rom[432] = 12'h000;
rom[433] = 12'h000;
rom[434] = 12'h00f;
rom[435] = 12'h00f;
rom[436] = 12'h00f;
rom[437] = 12'h00f;
rom[438] = 12'h00f;
rom[439] = 12'h00f;
rom[440] = 12'h000;
rom[441] = 12'h000;
rom[442] = 12'h000;
rom[443] = 12'h000;
rom[444] = 12'h007;
rom[445] = 12'h007;
rom[446] = 12'h000;
rom[447] = 12'h000;
rom[448] = 12'h007;
rom[449] = 12'h007;
rom[450] = 12'h000;
rom[451] = 12'h000;
rom[452] = 12'h000;
rom[453] = 12'h000;
rom[454] = 12'h000;
rom[455] = 12'h000;
rom[456] = 12'h000;
rom[457] = 12'h000;
rom[458] = 12'h000;
rom[459] = 12'h000;
rom[460] = 12'h00f;
rom[461] = 12'h00f;
rom[462] = 12'h00f;
rom[463] = 12'h00f;
rom[464] = 12'h00f;
rom[465] = 12'h00f;
rom[466] = 12'h000;
rom[467] = 12'h000;
rom[468] = 12'h000;
rom[469] = 12'h000;
rom[470] = 12'h000;
rom[471] = 12'h000;
rom[472] = 12'h007;
rom[473] = 12'h007;
rom[474] = 12'h000;
rom[475] = 12'h000;
rom[476] = 12'h000;
rom[477] = 12'h000;
rom[478] = 12'h000;
rom[479] = 12'h000;
rom[480] = 12'h000;
rom[481] = 12'h000;
rom[482] = 12'h000;
rom[483] = 12'h000;
rom[484] = 12'h000;
rom[485] = 12'h000;
rom[486] = 12'h000;
rom[487] = 12'h000;
rom[488] = 12'h00f;
rom[489] = 12'h00f;
rom[490] = 12'h00f;
rom[491] = 12'h00f;
rom[492] = 12'h000;
rom[493] = 12'h000;
rom[494] = 12'h000;
rom[495] = 12'h000;
rom[496] = 12'h000;
rom[497] = 12'h000;
rom[498] = 12'h007;
rom[499] = 12'h007;
rom[500] = 12'h000;
rom[501] = 12'h000;
rom[502] = 12'h000;
rom[503] = 12'h000;
rom[504] = 12'h000;
rom[505] = 12'h000;
rom[506] = 12'h000;
rom[507] = 12'h000;
rom[508] = 12'h000;
rom[509] = 12'h000;
rom[510] = 12'h000;
rom[511] = 12'h000;
rom[512] = 12'h000;
rom[513] = 12'h000;
rom[514] = 12'h00f;
rom[515] = 12'h00f;
rom[516] = 12'h00f;
rom[517] = 12'h00f;
rom[518] = 12'h000;
rom[519] = 12'h000;
rom[520] = 12'h000;
rom[521] = 12'h000;
rom[522] = 12'h007;
rom[523] = 12'h007;
rom[524] = 12'h000;
rom[525] = 12'h000;
rom[526] = 12'h000;
rom[527] = 12'h000;
rom[528] = 12'h007;
rom[529] = 12'h007;
rom[530] = 12'h000;
rom[531] = 12'h000;
rom[532] = 12'h007;
rom[533] = 12'h007;
rom[534] = 12'h000;
rom[535] = 12'h000;
rom[536] = 12'h007;
rom[537] = 12'h007;
rom[538] = 12'h000;
rom[539] = 12'h000;
rom[540] = 12'h000;
rom[541] = 12'h000;
rom[542] = 12'h00f;
rom[543] = 12'h00f;
rom[544] = 12'h000;
rom[545] = 12'h000;
rom[546] = 12'h000;
rom[547] = 12'h000;
rom[548] = 12'h007;
rom[549] = 12'h007;
rom[550] = 12'h000;
rom[551] = 12'h000;
rom[552] = 12'h000;
rom[553] = 12'h000;
rom[554] = 12'h007;
rom[555] = 12'h007;
rom[556] = 12'h000;
rom[557] = 12'h000;
rom[558] = 12'h007;
rom[559] = 12'h007;
rom[560] = 12'h000;
rom[561] = 12'h000;
rom[562] = 12'h007;
rom[563] = 12'h007;
rom[564] = 12'h000;
rom[565] = 12'h000;
rom[566] = 12'h000;
rom[567] = 12'h000;
rom[568] = 12'h00f;
rom[569] = 12'h00f;
rom[570] = 12'h000;
rom[571] = 12'h000;
rom[572] = 12'h000;
rom[573] = 12'h000;
rom[574] = 12'h000;
rom[575] = 12'h000;
rom[576] = 12'h000;
rom[577] = 12'h000;
rom[578] = 12'h007;
rom[579] = 12'h007;
rom[580] = 12'h000;
rom[581] = 12'h000;
rom[582] = 12'h007;
rom[583] = 12'h007;
rom[584] = 12'h000;
rom[585] = 12'h000;
rom[586] = 12'h007;
rom[587] = 12'h007;
rom[588] = 12'h000;
rom[589] = 12'h000;
rom[590] = 12'h007;
rom[591] = 12'h007;
rom[592] = 12'h000;
rom[593] = 12'h000;
rom[594] = 12'h000;
rom[595] = 12'h000;
rom[596] = 12'h000;
rom[597] = 12'h000;
rom[598] = 12'h000;
rom[599] = 12'h000;
rom[600] = 12'h000;
rom[601] = 12'h000;
rom[602] = 12'h000;
rom[603] = 12'h000;
rom[604] = 12'h007;
rom[605] = 12'h007;
rom[606] = 12'h000;
rom[607] = 12'h000;
rom[608] = 12'h007;
rom[609] = 12'h007;
rom[610] = 12'h000;
rom[611] = 12'h000;
rom[612] = 12'h007;
rom[613] = 12'h007;
rom[614] = 12'h000;
rom[615] = 12'h000;
rom[616] = 12'h007;
rom[617] = 12'h007;
rom[618] = 12'h000;
rom[619] = 12'h000;
rom[620] = 12'h000;
rom[621] = 12'h000;
rom[622] = 12'h000;
rom[623] = 12'h000;
rom[624] = 12'h000;
rom[625] = 12'h000;
rom[626] = 12'h007;
rom[627] = 12'h007;
rom[628] = 12'h000;
rom[629] = 12'h000;
rom[630] = 12'h000;
rom[631] = 12'h000;
rom[632] = 12'h007;
rom[633] = 12'h007;
rom[634] = 12'h000;
rom[635] = 12'h000;
rom[636] = 12'h007;
rom[637] = 12'h007;
rom[638] = 12'h000;
rom[639] = 12'h000;
rom[640] = 12'h007;
rom[641] = 12'h007;
rom[642] = 12'h000;
rom[643] = 12'h000;
rom[644] = 12'h000;
rom[645] = 12'h000;
rom[646] = 12'h00f;
rom[647] = 12'h00f;
rom[648] = 12'h000;
rom[649] = 12'h000;
rom[650] = 12'h000;
rom[651] = 12'h000;
rom[652] = 12'h007;
rom[653] = 12'h007;
rom[654] = 12'h000;
rom[655] = 12'h000;
rom[656] = 12'h000;
rom[657] = 12'h000;
rom[658] = 12'h007;
rom[659] = 12'h007;
rom[660] = 12'h000;
rom[661] = 12'h000;
rom[662] = 12'h007;
rom[663] = 12'h007;
rom[664] = 12'h000;
rom[665] = 12'h000;
rom[666] = 12'h007;
rom[667] = 12'h007;
rom[668] = 12'h000;
rom[669] = 12'h000;
rom[670] = 12'h000;
rom[671] = 12'h000;
rom[672] = 12'h00f;
rom[673] = 12'h00f;
rom[674] = 12'h000;
rom[675] = 12'h000;
rom[676] = 12'h000;
rom[677] = 12'h000;
rom[678] = 12'h000;
rom[679] = 12'h000;
rom[680] = 12'h007;
rom[681] = 12'h007;
rom[682] = 12'h000;
rom[683] = 12'h000;
rom[684] = 12'h000;
rom[685] = 12'h000;
rom[686] = 12'h000;
rom[687] = 12'h000;
rom[688] = 12'h000;
rom[689] = 12'h000;
rom[690] = 12'h000;
rom[691] = 12'h000;
rom[692] = 12'h000;
rom[693] = 12'h000;
rom[694] = 12'h000;
rom[695] = 12'h000;
rom[696] = 12'h00f;
rom[697] = 12'h00f;
rom[698] = 12'h00f;
rom[699] = 12'h00f;
rom[700] = 12'h000;
rom[701] = 12'h000;
rom[702] = 12'h000;
rom[703] = 12'h000;
rom[704] = 12'h000;
rom[705] = 12'h000;
rom[706] = 12'h007;
rom[707] = 12'h007;
rom[708] = 12'h000;
rom[709] = 12'h000;
rom[710] = 12'h000;
rom[711] = 12'h000;
rom[712] = 12'h000;
rom[713] = 12'h000;
rom[714] = 12'h000;
rom[715] = 12'h000;
rom[716] = 12'h000;
rom[717] = 12'h000;
rom[718] = 12'h000;
rom[719] = 12'h000;
rom[720] = 12'h000;
rom[721] = 12'h000;
rom[722] = 12'h00f;
rom[723] = 12'h00f;
rom[724] = 12'h00f;
rom[725] = 12'h00f;
rom[726] = 12'h000;
rom[727] = 12'h000;
rom[728] = 12'h000;
rom[729] = 12'h000;
rom[730] = 12'h007;
rom[731] = 12'h007;
rom[732] = 12'h000;
rom[733] = 12'h000;
rom[734] = 12'h007;
rom[735] = 12'h007;
rom[736] = 12'h000;
rom[737] = 12'h000;
rom[738] = 12'h000;
rom[739] = 12'h000;
rom[740] = 12'h000;
rom[741] = 12'h000;
rom[742] = 12'h000;
rom[743] = 12'h000;
rom[744] = 12'h000;
rom[745] = 12'h000;
rom[746] = 12'h00f;
rom[747] = 12'h00f;
rom[748] = 12'h00f;
rom[749] = 12'h00f;
rom[750] = 12'h00f;
rom[751] = 12'h00f;
rom[752] = 12'h000;
rom[753] = 12'h000;
rom[754] = 12'h000;
rom[755] = 12'h000;
rom[756] = 12'h007;
rom[757] = 12'h007;
rom[758] = 12'h000;
rom[759] = 12'h000;
rom[760] = 12'h007;
rom[761] = 12'h007;
rom[762] = 12'h000;
rom[763] = 12'h000;
rom[764] = 12'h000;
rom[765] = 12'h000;
rom[766] = 12'h000;
rom[767] = 12'h000;
rom[768] = 12'h000;
rom[769] = 12'h000;
rom[770] = 12'h000;
rom[771] = 12'h000;
rom[772] = 12'h00f;
rom[773] = 12'h00f;
rom[774] = 12'h00f;
rom[775] = 12'h00f;
rom[776] = 12'h00f;
rom[777] = 12'h00f;
rom[778] = 12'h000;
rom[779] = 12'h000;
rom[780] = 12'h000;
rom[781] = 12'h000;
rom[782] = 12'h000;
rom[783] = 12'h000;
rom[784] = 12'h007;
rom[785] = 12'h007;
rom[786] = 12'h000;
rom[787] = 12'h000;
rom[788] = 12'h000;
rom[789] = 12'h000;
rom[790] = 12'h000;
rom[791] = 12'h000;
rom[792] = 12'h000;
rom[793] = 12'h000;
rom[794] = 12'h000;
rom[795] = 12'h000;
rom[796] = 12'h000;
rom[797] = 12'h000;
rom[798] = 12'h00f;
rom[799] = 12'h00f;
rom[800] = 12'h00f;
rom[801] = 12'h00f;
rom[802] = 12'h00f;
rom[803] = 12'h00f;
rom[804] = 12'h000;
rom[805] = 12'h000;
rom[806] = 12'h000;
rom[807] = 12'h000;
rom[808] = 12'h000;
rom[809] = 12'h000;
rom[810] = 12'h007;
rom[811] = 12'h007;
rom[812] = 12'h000;
rom[813] = 12'h000;
rom[814] = 12'h000;
rom[815] = 12'h000;
rom[816] = 12'h000;
rom[817] = 12'h000;
rom[818] = 12'h000;
rom[819] = 12'h000;
rom[820] = 12'h000;
rom[821] = 12'h000;
rom[822] = 12'h000;
rom[823] = 12'h000;
rom[824] = 12'h00f;
rom[825] = 12'h00f;
rom[826] = 12'h00f;
rom[827] = 12'h00f;
rom[828] = 12'h00f;
rom[829] = 12'h00f;
rom[830] = 12'h000;
rom[831] = 12'h000;
rom[832] = 12'h000;
rom[833] = 12'h000;
rom[834] = 12'h007;
rom[835] = 12'h007;
rom[836] = 12'h000;
rom[837] = 12'h000;
rom[838] = 12'h007;
rom[839] = 12'h007;
rom[840] = 12'h000;
rom[841] = 12'h000;
rom[842] = 12'h000;
rom[843] = 12'h000;
rom[844] = 12'h000;
rom[845] = 12'h000;
rom[846] = 12'h000;
rom[847] = 12'h000;
rom[848] = 12'h000;
rom[849] = 12'h000;
rom[850] = 12'h00f;
rom[851] = 12'h00f;
rom[852] = 12'h00f;
rom[853] = 12'h00f;
rom[854] = 12'h00f;
rom[855] = 12'h00f;
rom[856] = 12'h000;
rom[857] = 12'h000;
rom[858] = 12'h000;
rom[859] = 12'h000;
rom[860] = 12'h007;
rom[861] = 12'h007;
rom[862] = 12'h000;
rom[863] = 12'h000;
rom[864] = 12'h007;
rom[865] = 12'h007;
rom[866] = 12'h000;
rom[867] = 12'h000;
rom[868] = 12'h000;
rom[869] = 12'h000;
rom[870] = 12'h000;
rom[871] = 12'h000;
rom[872] = 12'h000;
rom[873] = 12'h000;
rom[874] = 12'h000;
rom[875] = 12'h000;
rom[876] = 12'h00f;
rom[877] = 12'h00f;
rom[878] = 12'h00f;
rom[879] = 12'h00f;
rom[880] = 12'h00f;
rom[881] = 12'h00f;
rom[882] = 12'h000;
rom[883] = 12'h000;
rom[884] = 12'h000;
rom[885] = 12'h000;
rom[886] = 12'h000;
rom[887] = 12'h000;
rom[888] = 12'h007;
rom[889] = 12'h007;
rom[890] = 12'h000;
rom[891] = 12'h000;
rom[892] = 12'h000;
rom[893] = 12'h000;
rom[894] = 12'h000;
rom[895] = 12'h000;
rom[896] = 12'h000;
rom[897] = 12'h000;
rom[898] = 12'h000;
rom[899] = 12'h000;
rom[900] = 12'h000;
rom[901] = 12'h000;
rom[902] = 12'h00f;
rom[903] = 12'h00f;
rom[904] = 12'h00f;
rom[905] = 12'h00f;
rom[906] = 12'h00f;
rom[907] = 12'h00f;
rom[908] = 12'h000;
rom[909] = 12'h000;
rom[910] = 12'h000;
rom[911] = 12'h000;
rom[912] = 12'h000;
rom[913] = 12'h000;
rom[914] = 12'h007;
rom[915] = 12'h007;
rom[916] = 12'h000;
rom[917] = 12'h000;
rom[918] = 12'h000;
rom[919] = 12'h000;
rom[920] = 12'h000;
rom[921] = 12'h000;
rom[922] = 12'h000;
rom[923] = 12'h000;
rom[924] = 12'h000;
rom[925] = 12'h000;
rom[926] = 12'h000;
rom[927] = 12'h000;
rom[928] = 12'h00f;
rom[929] = 12'h00f;
rom[930] = 12'h00f;
rom[931] = 12'h00f;
rom[932] = 12'h00f;
rom[933] = 12'h00f;
rom[934] = 12'h000;
rom[935] = 12'h000;
rom[936] = 12'h000;
rom[937] = 12'h000;
rom[938] = 12'h007;
rom[939] = 12'h007;
rom[940] = 12'h000;
rom[941] = 12'h000;
rom[942] = 12'h007;
rom[943] = 12'h007;
rom[944] = 12'h000;
rom[945] = 12'h000;
rom[946] = 12'h000;
rom[947] = 12'h000;
rom[948] = 12'h000;
rom[949] = 12'h000;
rom[950] = 12'h000;
rom[951] = 12'h000;
rom[952] = 12'h000;
rom[953] = 12'h000;
rom[954] = 12'h00f;
rom[955] = 12'h00f;
rom[956] = 12'h00f;
rom[957] = 12'h00f;
rom[958] = 12'h00f;
rom[959] = 12'h00f;
rom[960] = 12'h000;
rom[961] = 12'h000;
rom[962] = 12'h000;
rom[963] = 12'h000;
rom[964] = 12'h007;
rom[965] = 12'h007;
rom[966] = 12'h000;
rom[967] = 12'h000;
rom[968] = 12'h007;
rom[969] = 12'h007;
rom[970] = 12'h000;
rom[971] = 12'h000;
rom[972] = 12'h000;
rom[973] = 12'h000;
rom[974] = 12'h000;
rom[975] = 12'h000;
rom[976] = 12'h000;
rom[977] = 12'h000;
rom[978] = 12'h000;
rom[979] = 12'h000;
rom[980] = 12'h00f;
rom[981] = 12'h00f;
rom[982] = 12'h00f;
rom[983] = 12'h00f;
rom[984] = 12'h00f;
rom[985] = 12'h00f;
rom[986] = 12'h000;
rom[987] = 12'h000;
rom[988] = 12'h000;
rom[989] = 12'h000;
rom[990] = 12'h000;
rom[991] = 12'h000;
rom[992] = 12'h007;
rom[993] = 12'h007;
rom[994] = 12'h000;
rom[995] = 12'h000;
rom[996] = 12'h000;
rom[997] = 12'h000;
rom[998] = 12'h007;
rom[999] = 12'h007;
rom[1000] = 12'h000;
rom[1001] = 12'h000;
rom[1002] = 12'h007;
rom[1003] = 12'h007;
rom[1004] = 12'h000;
rom[1005] = 12'h000;
rom[1006] = 12'h000;
rom[1007] = 12'h000;
rom[1008] = 12'h00f;
rom[1009] = 12'h00f;
rom[1010] = 12'h00f;
rom[1011] = 12'h00f;
rom[1012] = 12'h000;
rom[1013] = 12'h000;
rom[1014] = 12'h000;
rom[1015] = 12'h000;
rom[1016] = 12'h000;
rom[1017] = 12'h000;
rom[1018] = 12'h007;
rom[1019] = 12'h007;
rom[1020] = 12'h000;
rom[1021] = 12'h000;
rom[1022] = 12'h000;
rom[1023] = 12'h000;
rom[1024] = 12'h007;
rom[1025] = 12'h007;
rom[1026] = 12'h000;
rom[1027] = 12'h000;
rom[1028] = 12'h007;
rom[1029] = 12'h007;
rom[1030] = 12'h000;
rom[1031] = 12'h000;
rom[1032] = 12'h000;
rom[1033] = 12'h000;
rom[1034] = 12'h00f;
rom[1035] = 12'h00f;
rom[1036] = 12'h00f;
rom[1037] = 12'h00f;
rom[1038] = 12'h000;
rom[1039] = 12'h000;
rom[1040] = 12'h000;
rom[1041] = 12'h000;
rom[1042] = 12'h007;
rom[1043] = 12'h007;
rom[1044] = 12'h000;
rom[1045] = 12'h000;
rom[1046] = 12'h000;
rom[1047] = 12'h000;
rom[1048] = 12'h007;
rom[1049] = 12'h007;
rom[1050] = 12'h000;
rom[1051] = 12'h000;
rom[1052] = 12'h007;
rom[1053] = 12'h007;
rom[1054] = 12'h000;
rom[1055] = 12'h000;
rom[1056] = 12'h007;
rom[1057] = 12'h007;
rom[1058] = 12'h000;
rom[1059] = 12'h000;
rom[1060] = 12'h000;
rom[1061] = 12'h000;
rom[1062] = 12'h00f;
rom[1063] = 12'h00f;
rom[1064] = 12'h000;
rom[1065] = 12'h000;
rom[1066] = 12'h000;
rom[1067] = 12'h000;
rom[1068] = 12'h007;
rom[1069] = 12'h007;
rom[1070] = 12'h000;
rom[1071] = 12'h000;
rom[1072] = 12'h000;
rom[1073] = 12'h000;
rom[1074] = 12'h007;
rom[1075] = 12'h007;
rom[1076] = 12'h000;
rom[1077] = 12'h000;
rom[1078] = 12'h007;
rom[1079] = 12'h007;
rom[1080] = 12'h000;
rom[1081] = 12'h000;
rom[1082] = 12'h007;
rom[1083] = 12'h007;
rom[1084] = 12'h000;
rom[1085] = 12'h000;
rom[1086] = 12'h000;
rom[1087] = 12'h000;
rom[1088] = 12'h00f;
rom[1089] = 12'h00f;
rom[1090] = 12'h000;
rom[1091] = 12'h000;
rom[1092] = 12'h000;
rom[1093] = 12'h000;
rom[1094] = 12'h000;
rom[1095] = 12'h000;
rom[1096] = 12'h000;
rom[1097] = 12'h000;
rom[1098] = 12'h007;
rom[1099] = 12'h007;
rom[1100] = 12'h000;
rom[1101] = 12'h000;
rom[1102] = 12'h007;
rom[1103] = 12'h007;
rom[1104] = 12'h000;
rom[1105] = 12'h000;
rom[1106] = 12'h007;
rom[1107] = 12'h007;
rom[1108] = 12'h000;
rom[1109] = 12'h000;
rom[1110] = 12'h007;
rom[1111] = 12'h007;
rom[1112] = 12'h000;
rom[1113] = 12'h000;
rom[1114] = 12'h000;
rom[1115] = 12'h000;
rom[1116] = 12'h000;
rom[1117] = 12'h000;
rom[1118] = 12'h000;
rom[1119] = 12'h000;
rom[1120] = 12'h000;
rom[1121] = 12'h000;
rom[1122] = 12'h000;
rom[1123] = 12'h000;
rom[1124] = 12'h007;
rom[1125] = 12'h007;
rom[1126] = 12'h000;
rom[1127] = 12'h000;
rom[1128] = 12'h007;
rom[1129] = 12'h007;
rom[1130] = 12'h000;
rom[1131] = 12'h000;
rom[1132] = 12'h007;
rom[1133] = 12'h007;
rom[1134] = 12'h000;
rom[1135] = 12'h000;
rom[1136] = 12'h007;
rom[1137] = 12'h007;
rom[1138] = 12'h000;
rom[1139] = 12'h000;
rom[1140] = 12'h000;
rom[1141] = 12'h000;
rom[1142] = 12'h000;
rom[1143] = 12'h000;
rom[1144] = 12'h000;
rom[1145] = 12'h000;
rom[1146] = 12'h000;
rom[1147] = 12'h000;
rom[1148] = 12'h000;
rom[1149] = 12'h000;
rom[1150] = 12'h000;
rom[1151] = 12'h000;
rom[1152] = 12'h000;
rom[1153] = 12'h000;
rom[1154] = 12'h000;
rom[1155] = 12'h000;
rom[1156] = 12'h000;
rom[1157] = 12'h000;
rom[1158] = 12'h000;
rom[1159] = 12'h000;
rom[1160] = 12'h000;
rom[1161] = 12'h000;
rom[1162] = 12'h000;
rom[1163] = 12'h000;
rom[1164] = 12'h000;
rom[1165] = 12'h000;
rom[1166] = 12'h000;
rom[1167] = 12'h000;
rom[1168] = 12'h000;
rom[1169] = 12'h000;
rom[1170] = 12'h000;
rom[1171] = 12'h000;
rom[1172] = 12'h000;
rom[1173] = 12'h000;
rom[1174] = 12'h000;
rom[1175] = 12'h000;
rom[1176] = 12'h000;
rom[1177] = 12'h000;
rom[1178] = 12'h000;
rom[1179] = 12'h000;
rom[1180] = 12'h000;
rom[1181] = 12'h000;
rom[1182] = 12'h000;
rom[1183] = 12'h000;
rom[1184] = 12'h000;
rom[1185] = 12'h000;
rom[1186] = 12'h000;
rom[1187] = 12'h000;
rom[1188] = 12'h000;
rom[1189] = 12'h000;
rom[1190] = 12'h000;
rom[1191] = 12'h000;
rom[1192] = 12'h000;
rom[1193] = 12'h000;
rom[1194] = 12'h000;
rom[1195] = 12'h000;
  end
  endmodule

    module dash_rom (                       //два
  input  wire    [13:0]     addr,
  output wire    [11:0]     word
);

  logic [11:0] rom [(46 * 26)];

  assign word = rom[addr];

  initial begin
rom[0] = 12'h000;
rom[1] = 12'h000;
rom[2] = 12'h000;
rom[3] = 12'h000;
rom[4] = 12'h000;
rom[5] = 12'h000;
rom[6] = 12'h000;
rom[7] = 12'h000;
rom[8] = 12'h000;
rom[9] = 12'h000;
rom[10] = 12'h000;
rom[11] = 12'h000;
rom[12] = 12'h000;
rom[13] = 12'h000;
rom[14] = 12'h000;
rom[15] = 12'h000;
rom[16] = 12'h000;
rom[17] = 12'h000;
rom[18] = 12'h000;
rom[19] = 12'h000;
rom[20] = 12'h000;
rom[21] = 12'h000;
rom[22] = 12'h000;
rom[23] = 12'h000;
rom[24] = 12'h000;
rom[25] = 12'h000;
rom[26] = 12'h000;
rom[27] = 12'h000;
rom[28] = 12'h000;
rom[29] = 12'h000;
rom[30] = 12'h000;
rom[31] = 12'h000;
rom[32] = 12'h000;
rom[33] = 12'h000;
rom[34] = 12'h000;
rom[35] = 12'h000;
rom[36] = 12'h000;
rom[37] = 12'h000;
rom[38] = 12'h000;
rom[39] = 12'h000;
rom[40] = 12'h000;
rom[41] = 12'h000;
rom[42] = 12'h000;
rom[43] = 12'h000;
rom[44] = 12'h000;
rom[45] = 12'h000;
rom[46] = 12'h000;
rom[47] = 12'h000;
rom[48] = 12'h000;
rom[49] = 12'h000;
rom[50] = 12'h000;
rom[51] = 12'h000;
rom[52] = 12'h000;
rom[53] = 12'h000;
rom[54] = 12'h000;
rom[55] = 12'h000;
rom[56] = 12'h00f;
rom[57] = 12'h00f;
rom[58] = 12'h00f;
rom[59] = 12'h00f;
rom[60] = 12'h00f;
rom[61] = 12'h00f;
rom[62] = 12'h00f;
rom[63] = 12'h00f;
rom[64] = 12'h00f;
rom[65] = 12'h00f;
rom[66] = 12'h00f;
rom[67] = 12'h00f;
rom[68] = 12'h00f;
rom[69] = 12'h00f;
rom[70] = 12'h00f;
rom[71] = 12'h00f;
rom[72] = 12'h00f;
rom[73] = 12'h00f;
rom[74] = 12'h000;
rom[75] = 12'h000;
rom[76] = 12'h000;
rom[77] = 12'h000;
rom[78] = 12'h000;
rom[79] = 12'h000;
rom[80] = 12'h000;
rom[81] = 12'h000;
rom[82] = 12'h00f;
rom[83] = 12'h00f;
rom[84] = 12'h00f;
rom[85] = 12'h00f;
rom[86] = 12'h00f;
rom[87] = 12'h00f;
rom[88] = 12'h00f;
rom[89] = 12'h00f;
rom[90] = 12'h00f;
rom[91] = 12'h00f;
rom[92] = 12'h00f;
rom[93] = 12'h00f;
rom[94] = 12'h00f;
rom[95] = 12'h00f;
rom[96] = 12'h00f;
rom[97] = 12'h00f;
rom[98] = 12'h00f;
rom[99] = 12'h00f;
rom[100] = 12'h000;
rom[101] = 12'h000;
rom[102] = 12'h000;
rom[103] = 12'h000;
rom[104] = 12'h000;
rom[105] = 12'h000;
rom[106] = 12'h007;
rom[107] = 12'h007;
rom[108] = 12'h000;
rom[109] = 12'h000;
rom[110] = 12'h00f;
rom[111] = 12'h00f;
rom[112] = 12'h00f;
rom[113] = 12'h00f;
rom[114] = 12'h00f;
rom[115] = 12'h00f;
rom[116] = 12'h00f;
rom[117] = 12'h00f;
rom[118] = 12'h00f;
rom[119] = 12'h00f;
rom[120] = 12'h00f;
rom[121] = 12'h00f;
rom[122] = 12'h00f;
rom[123] = 12'h00f;
rom[124] = 12'h000;
rom[125] = 12'h000;
rom[126] = 12'h00f;
rom[127] = 12'h00f;
rom[128] = 12'h000;
rom[129] = 12'h000;
rom[130] = 12'h000;
rom[131] = 12'h000;
rom[132] = 12'h007;
rom[133] = 12'h007;
rom[134] = 12'h000;
rom[135] = 12'h000;
rom[136] = 12'h00f;
rom[137] = 12'h00f;
rom[138] = 12'h00f;
rom[139] = 12'h00f;
rom[140] = 12'h00f;
rom[141] = 12'h00f;
rom[142] = 12'h00f;
rom[143] = 12'h00f;
rom[144] = 12'h00f;
rom[145] = 12'h00f;
rom[146] = 12'h00f;
rom[147] = 12'h00f;
rom[148] = 12'h00f;
rom[149] = 12'h00f;
rom[150] = 12'h000;
rom[151] = 12'h000;
rom[152] = 12'h00f;
rom[153] = 12'h00f;
rom[154] = 12'h000;
rom[155] = 12'h000;
rom[156] = 12'h000;
rom[157] = 12'h000;
rom[158] = 12'h000;
rom[159] = 12'h000;
rom[160] = 12'h007;
rom[161] = 12'h007;
rom[162] = 12'h000;
rom[163] = 12'h000;
rom[164] = 12'h00f;
rom[165] = 12'h00f;
rom[166] = 12'h00f;
rom[167] = 12'h00f;
rom[168] = 12'h00f;
rom[169] = 12'h00f;
rom[170] = 12'h00f;
rom[171] = 12'h00f;
rom[172] = 12'h00f;
rom[173] = 12'h00f;
rom[174] = 12'h000;
rom[175] = 12'h000;
rom[176] = 12'h00f;
rom[177] = 12'h00f;
rom[178] = 12'h00f;
rom[179] = 12'h00f;
rom[180] = 12'h000;
rom[181] = 12'h000;
rom[182] = 12'h000;
rom[183] = 12'h000;
rom[184] = 12'h000;
rom[185] = 12'h000;
rom[186] = 12'h007;
rom[187] = 12'h007;
rom[188] = 12'h000;
rom[189] = 12'h000;
rom[190] = 12'h00f;
rom[191] = 12'h00f;
rom[192] = 12'h00f;
rom[193] = 12'h00f;
rom[194] = 12'h00f;
rom[195] = 12'h00f;
rom[196] = 12'h00f;
rom[197] = 12'h00f;
rom[198] = 12'h00f;
rom[199] = 12'h00f;
rom[200] = 12'h000;
rom[201] = 12'h000;
rom[202] = 12'h00f;
rom[203] = 12'h00f;
rom[204] = 12'h00f;
rom[205] = 12'h00f;
rom[206] = 12'h000;
rom[207] = 12'h000;
rom[208] = 12'h000;
rom[209] = 12'h000;
rom[210] = 12'h007;
rom[211] = 12'h007;
rom[212] = 12'h000;
rom[213] = 12'h000;
rom[214] = 12'h007;
rom[215] = 12'h007;
rom[216] = 12'h000;
rom[217] = 12'h000;
rom[218] = 12'h000;
rom[219] = 12'h000;
rom[220] = 12'h000;
rom[221] = 12'h000;
rom[222] = 12'h000;
rom[223] = 12'h000;
rom[224] = 12'h000;
rom[225] = 12'h000;
rom[226] = 12'h00f;
rom[227] = 12'h00f;
rom[228] = 12'h00f;
rom[229] = 12'h00f;
rom[230] = 12'h00f;
rom[231] = 12'h00f;
rom[232] = 12'h000;
rom[233] = 12'h000;
rom[234] = 12'h000;
rom[235] = 12'h000;
rom[236] = 12'h007;
rom[237] = 12'h007;
rom[238] = 12'h000;
rom[239] = 12'h000;
rom[240] = 12'h007;
rom[241] = 12'h007;
rom[242] = 12'h000;
rom[243] = 12'h000;
rom[244] = 12'h000;
rom[245] = 12'h000;
rom[246] = 12'h000;
rom[247] = 12'h000;
rom[248] = 12'h000;
rom[249] = 12'h000;
rom[250] = 12'h000;
rom[251] = 12'h000;
rom[252] = 12'h00f;
rom[253] = 12'h00f;
rom[254] = 12'h00f;
rom[255] = 12'h00f;
rom[256] = 12'h00f;
rom[257] = 12'h00f;
rom[258] = 12'h000;
rom[259] = 12'h000;
rom[260] = 12'h000;
rom[261] = 12'h000;
rom[262] = 12'h000;
rom[263] = 12'h000;
rom[264] = 12'h007;
rom[265] = 12'h007;
rom[266] = 12'h000;
rom[267] = 12'h000;
rom[268] = 12'h000;
rom[269] = 12'h000;
rom[270] = 12'h000;
rom[271] = 12'h000;
rom[272] = 12'h000;
rom[273] = 12'h000;
rom[274] = 12'h000;
rom[275] = 12'h000;
rom[276] = 12'h000;
rom[277] = 12'h000;
rom[278] = 12'h00f;
rom[279] = 12'h00f;
rom[280] = 12'h00f;
rom[281] = 12'h00f;
rom[282] = 12'h00f;
rom[283] = 12'h00f;
rom[284] = 12'h000;
rom[285] = 12'h000;
rom[286] = 12'h000;
rom[287] = 12'h000;
rom[288] = 12'h000;
rom[289] = 12'h000;
rom[290] = 12'h007;
rom[291] = 12'h007;
rom[292] = 12'h000;
rom[293] = 12'h000;
rom[294] = 12'h000;
rom[295] = 12'h000;
rom[296] = 12'h000;
rom[297] = 12'h000;
rom[298] = 12'h000;
rom[299] = 12'h000;
rom[300] = 12'h000;
rom[301] = 12'h000;
rom[302] = 12'h000;
rom[303] = 12'h000;
rom[304] = 12'h00f;
rom[305] = 12'h00f;
rom[306] = 12'h00f;
rom[307] = 12'h00f;
rom[308] = 12'h00f;
rom[309] = 12'h00f;
rom[310] = 12'h000;
rom[311] = 12'h000;
rom[312] = 12'h000;
rom[313] = 12'h000;
rom[314] = 12'h007;
rom[315] = 12'h007;
rom[316] = 12'h000;
rom[317] = 12'h000;
rom[318] = 12'h007;
rom[319] = 12'h007;
rom[320] = 12'h000;
rom[321] = 12'h000;
rom[322] = 12'h000;
rom[323] = 12'h000;
rom[324] = 12'h000;
rom[325] = 12'h000;
rom[326] = 12'h000;
rom[327] = 12'h000;
rom[328] = 12'h000;
rom[329] = 12'h000;
rom[330] = 12'h00f;
rom[331] = 12'h00f;
rom[332] = 12'h00f;
rom[333] = 12'h00f;
rom[334] = 12'h00f;
rom[335] = 12'h00f;
rom[336] = 12'h000;
rom[337] = 12'h000;
rom[338] = 12'h000;
rom[339] = 12'h000;
rom[340] = 12'h007;
rom[341] = 12'h007;
rom[342] = 12'h000;
rom[343] = 12'h000;
rom[344] = 12'h007;
rom[345] = 12'h007;
rom[346] = 12'h000;
rom[347] = 12'h000;
rom[348] = 12'h000;
rom[349] = 12'h000;
rom[350] = 12'h000;
rom[351] = 12'h000;
rom[352] = 12'h000;
rom[353] = 12'h000;
rom[354] = 12'h000;
rom[355] = 12'h000;
rom[356] = 12'h00f;
rom[357] = 12'h00f;
rom[358] = 12'h00f;
rom[359] = 12'h00f;
rom[360] = 12'h00f;
rom[361] = 12'h00f;
rom[362] = 12'h000;
rom[363] = 12'h000;
rom[364] = 12'h000;
rom[365] = 12'h000;
rom[366] = 12'h000;
rom[367] = 12'h000;
rom[368] = 12'h007;
rom[369] = 12'h007;
rom[370] = 12'h000;
rom[371] = 12'h000;
rom[372] = 12'h000;
rom[373] = 12'h000;
rom[374] = 12'h000;
rom[375] = 12'h000;
rom[376] = 12'h000;
rom[377] = 12'h000;
rom[378] = 12'h000;
rom[379] = 12'h000;
rom[380] = 12'h000;
rom[381] = 12'h000;
rom[382] = 12'h00f;
rom[383] = 12'h00f;
rom[384] = 12'h00f;
rom[385] = 12'h00f;
rom[386] = 12'h00f;
rom[387] = 12'h00f;
rom[388] = 12'h000;
rom[389] = 12'h000;
rom[390] = 12'h000;
rom[391] = 12'h000;
rom[392] = 12'h000;
rom[393] = 12'h000;
rom[394] = 12'h007;
rom[395] = 12'h007;
rom[396] = 12'h000;
rom[397] = 12'h000;
rom[398] = 12'h000;
rom[399] = 12'h000;
rom[400] = 12'h000;
rom[401] = 12'h000;
rom[402] = 12'h000;
rom[403] = 12'h000;
rom[404] = 12'h000;
rom[405] = 12'h000;
rom[406] = 12'h000;
rom[407] = 12'h000;
rom[408] = 12'h00f;
rom[409] = 12'h00f;
rom[410] = 12'h00f;
rom[411] = 12'h00f;
rom[412] = 12'h00f;
rom[413] = 12'h00f;
rom[414] = 12'h000;
rom[415] = 12'h000;
rom[416] = 12'h000;
rom[417] = 12'h000;
rom[418] = 12'h007;
rom[419] = 12'h007;
rom[420] = 12'h000;
rom[421] = 12'h000;
rom[422] = 12'h007;
rom[423] = 12'h007;
rom[424] = 12'h000;
rom[425] = 12'h000;
rom[426] = 12'h000;
rom[427] = 12'h000;
rom[428] = 12'h000;
rom[429] = 12'h000;
rom[430] = 12'h000;
rom[431] = 12'h000;
rom[432] = 12'h000;
rom[433] = 12'h000;
rom[434] = 12'h00f;
rom[435] = 12'h00f;
rom[436] = 12'h00f;
rom[437] = 12'h00f;
rom[438] = 12'h00f;
rom[439] = 12'h00f;
rom[440] = 12'h000;
rom[441] = 12'h000;
rom[442] = 12'h000;
rom[443] = 12'h000;
rom[444] = 12'h007;
rom[445] = 12'h007;
rom[446] = 12'h000;
rom[447] = 12'h000;
rom[448] = 12'h007;
rom[449] = 12'h007;
rom[450] = 12'h000;
rom[451] = 12'h000;
rom[452] = 12'h000;
rom[453] = 12'h000;
rom[454] = 12'h000;
rom[455] = 12'h000;
rom[456] = 12'h000;
rom[457] = 12'h000;
rom[458] = 12'h000;
rom[459] = 12'h000;
rom[460] = 12'h00f;
rom[461] = 12'h00f;
rom[462] = 12'h00f;
rom[463] = 12'h00f;
rom[464] = 12'h00f;
rom[465] = 12'h00f;
rom[466] = 12'h000;
rom[467] = 12'h000;
rom[468] = 12'h000;
rom[469] = 12'h000;
rom[470] = 12'h000;
rom[471] = 12'h000;
rom[472] = 12'h007;
rom[473] = 12'h007;
rom[474] = 12'h000;
rom[475] = 12'h000;
rom[476] = 12'h000;
rom[477] = 12'h000;
rom[478] = 12'h000;
rom[479] = 12'h000;
rom[480] = 12'h000;
rom[481] = 12'h000;
rom[482] = 12'h000;
rom[483] = 12'h000;
rom[484] = 12'h000;
rom[485] = 12'h000;
rom[486] = 12'h000;
rom[487] = 12'h000;
rom[488] = 12'h00f;
rom[489] = 12'h00f;
rom[490] = 12'h00f;
rom[491] = 12'h00f;
rom[492] = 12'h000;
rom[493] = 12'h000;
rom[494] = 12'h000;
rom[495] = 12'h000;
rom[496] = 12'h000;
rom[497] = 12'h000;
rom[498] = 12'h007;
rom[499] = 12'h007;
rom[500] = 12'h000;
rom[501] = 12'h000;
rom[502] = 12'h000;
rom[503] = 12'h000;
rom[504] = 12'h000;
rom[505] = 12'h000;
rom[506] = 12'h000;
rom[507] = 12'h000;
rom[508] = 12'h000;
rom[509] = 12'h000;
rom[510] = 12'h000;
rom[511] = 12'h000;
rom[512] = 12'h000;
rom[513] = 12'h000;
rom[514] = 12'h00f;
rom[515] = 12'h00f;
rom[516] = 12'h00f;
rom[517] = 12'h00f;
rom[518] = 12'h000;
rom[519] = 12'h000;
rom[520] = 12'h000;
rom[521] = 12'h000;
rom[522] = 12'h007;
rom[523] = 12'h007;
rom[524] = 12'h000;
rom[525] = 12'h000;
rom[526] = 12'h00f;
rom[527] = 12'h00f;
rom[528] = 12'h00f;
rom[529] = 12'h00f;
rom[530] = 12'h00f;
rom[531] = 12'h00f;
rom[532] = 12'h00f;
rom[533] = 12'h00f;
rom[534] = 12'h00f;
rom[535] = 12'h00f;
rom[536] = 12'h00f;
rom[537] = 12'h00f;
rom[538] = 12'h00f;
rom[539] = 12'h00f;
rom[540] = 12'h000;
rom[541] = 12'h000;
rom[542] = 12'h00f;
rom[543] = 12'h00f;
rom[544] = 12'h000;
rom[545] = 12'h000;
rom[546] = 12'h000;
rom[547] = 12'h000;
rom[548] = 12'h007;
rom[549] = 12'h007;
rom[550] = 12'h000;
rom[551] = 12'h000;
rom[552] = 12'h00f;
rom[553] = 12'h00f;
rom[554] = 12'h00f;
rom[555] = 12'h00f;
rom[556] = 12'h00f;
rom[557] = 12'h00f;
rom[558] = 12'h00f;
rom[559] = 12'h00f;
rom[560] = 12'h00f;
rom[561] = 12'h00f;
rom[562] = 12'h00f;
rom[563] = 12'h00f;
rom[564] = 12'h00f;
rom[565] = 12'h00f;
rom[566] = 12'h000;
rom[567] = 12'h000;
rom[568] = 12'h00f;
rom[569] = 12'h00f;
rom[570] = 12'h000;
rom[571] = 12'h000;
rom[572] = 12'h000;
rom[573] = 12'h000;
rom[574] = 12'h000;
rom[575] = 12'h000;
rom[576] = 12'h00f;
rom[577] = 12'h00f;
rom[578] = 12'h00f;
rom[579] = 12'h00f;
rom[580] = 12'h00f;
rom[581] = 12'h00f;
rom[582] = 12'h00f;
rom[583] = 12'h00f;
rom[584] = 12'h00f;
rom[585] = 12'h00f;
rom[586] = 12'h00f;
rom[587] = 12'h00f;
rom[588] = 12'h00f;
rom[589] = 12'h00f;
rom[590] = 12'h00f;
rom[591] = 12'h00f;
rom[592] = 12'h00f;
rom[593] = 12'h00f;
rom[594] = 12'h000;
rom[595] = 12'h000;
rom[596] = 12'h000;
rom[597] = 12'h000;
rom[598] = 12'h000;
rom[599] = 12'h000;
rom[600] = 12'h000;
rom[601] = 12'h000;
rom[602] = 12'h00f;
rom[603] = 12'h00f;
rom[604] = 12'h00f;
rom[605] = 12'h00f;
rom[606] = 12'h00f;
rom[607] = 12'h00f;
rom[608] = 12'h00f;
rom[609] = 12'h00f;
rom[610] = 12'h00f;
rom[611] = 12'h00f;
rom[612] = 12'h00f;
rom[613] = 12'h00f;
rom[614] = 12'h00f;
rom[615] = 12'h00f;
rom[616] = 12'h00f;
rom[617] = 12'h00f;
rom[618] = 12'h00f;
rom[619] = 12'h00f;
rom[620] = 12'h000;
rom[621] = 12'h000;
rom[622] = 12'h000;
rom[623] = 12'h000;
rom[624] = 12'h000;
rom[625] = 12'h000;
rom[626] = 12'h00f;
rom[627] = 12'h00f;
rom[628] = 12'h000;
rom[629] = 12'h000;
rom[630] = 12'h00f;
rom[631] = 12'h00f;
rom[632] = 12'h00f;
rom[633] = 12'h00f;
rom[634] = 12'h00f;
rom[635] = 12'h00f;
rom[636] = 12'h00f;
rom[637] = 12'h00f;
rom[638] = 12'h00f;
rom[639] = 12'h00f;
rom[640] = 12'h00f;
rom[641] = 12'h00f;
rom[642] = 12'h00f;
rom[643] = 12'h00f;
rom[644] = 12'h000;
rom[645] = 12'h000;
rom[646] = 12'h007;
rom[647] = 12'h007;
rom[648] = 12'h000;
rom[649] = 12'h000;
rom[650] = 12'h000;
rom[651] = 12'h000;
rom[652] = 12'h00f;
rom[653] = 12'h00f;
rom[654] = 12'h000;
rom[655] = 12'h000;
rom[656] = 12'h00f;
rom[657] = 12'h00f;
rom[658] = 12'h00f;
rom[659] = 12'h00f;
rom[660] = 12'h00f;
rom[661] = 12'h00f;
rom[662] = 12'h00f;
rom[663] = 12'h00f;
rom[664] = 12'h00f;
rom[665] = 12'h00f;
rom[666] = 12'h00f;
rom[667] = 12'h00f;
rom[668] = 12'h00f;
rom[669] = 12'h00f;
rom[670] = 12'h000;
rom[671] = 12'h000;
rom[672] = 12'h007;
rom[673] = 12'h007;
rom[674] = 12'h000;
rom[675] = 12'h000;
rom[676] = 12'h000;
rom[677] = 12'h000;
rom[678] = 12'h00f;
rom[679] = 12'h00f;
rom[680] = 12'h00f;
rom[681] = 12'h00f;
rom[682] = 12'h000;
rom[683] = 12'h000;
rom[684] = 12'h000;
rom[685] = 12'h000;
rom[686] = 12'h000;
rom[687] = 12'h000;
rom[688] = 12'h000;
rom[689] = 12'h000;
rom[690] = 12'h000;
rom[691] = 12'h000;
rom[692] = 12'h000;
rom[693] = 12'h000;
rom[694] = 12'h000;
rom[695] = 12'h000;
rom[696] = 12'h007;
rom[697] = 12'h007;
rom[698] = 12'h000;
rom[699] = 12'h000;
rom[700] = 12'h000;
rom[701] = 12'h000;
rom[702] = 12'h000;
rom[703] = 12'h000;
rom[704] = 12'h00f;
rom[705] = 12'h00f;
rom[706] = 12'h00f;
rom[707] = 12'h00f;
rom[708] = 12'h000;
rom[709] = 12'h000;
rom[710] = 12'h000;
rom[711] = 12'h000;
rom[712] = 12'h000;
rom[713] = 12'h000;
rom[714] = 12'h000;
rom[715] = 12'h000;
rom[716] = 12'h000;
rom[717] = 12'h000;
rom[718] = 12'h000;
rom[719] = 12'h000;
rom[720] = 12'h000;
rom[721] = 12'h000;
rom[722] = 12'h007;
rom[723] = 12'h007;
rom[724] = 12'h000;
rom[725] = 12'h000;
rom[726] = 12'h000;
rom[727] = 12'h000;
rom[728] = 12'h000;
rom[729] = 12'h000;
rom[730] = 12'h00f;
rom[731] = 12'h00f;
rom[732] = 12'h00f;
rom[733] = 12'h00f;
rom[734] = 12'h00f;
rom[735] = 12'h00f;
rom[736] = 12'h000;
rom[737] = 12'h000;
rom[738] = 12'h000;
rom[739] = 12'h000;
rom[740] = 12'h000;
rom[741] = 12'h000;
rom[742] = 12'h000;
rom[743] = 12'h000;
rom[744] = 12'h000;
rom[745] = 12'h000;
rom[746] = 12'h007;
rom[747] = 12'h007;
rom[748] = 12'h000;
rom[749] = 12'h000;
rom[750] = 12'h007;
rom[751] = 12'h007;
rom[752] = 12'h000;
rom[753] = 12'h000;
rom[754] = 12'h000;
rom[755] = 12'h000;
rom[756] = 12'h00f;
rom[757] = 12'h00f;
rom[758] = 12'h00f;
rom[759] = 12'h00f;
rom[760] = 12'h00f;
rom[761] = 12'h00f;
rom[762] = 12'h000;
rom[763] = 12'h000;
rom[764] = 12'h000;
rom[765] = 12'h000;
rom[766] = 12'h000;
rom[767] = 12'h000;
rom[768] = 12'h000;
rom[769] = 12'h000;
rom[770] = 12'h000;
rom[771] = 12'h000;
rom[772] = 12'h007;
rom[773] = 12'h007;
rom[774] = 12'h000;
rom[775] = 12'h000;
rom[776] = 12'h007;
rom[777] = 12'h007;
rom[778] = 12'h000;
rom[779] = 12'h000;
rom[780] = 12'h000;
rom[781] = 12'h000;
rom[782] = 12'h00f;
rom[783] = 12'h00f;
rom[784] = 12'h00f;
rom[785] = 12'h00f;
rom[786] = 12'h00f;
rom[787] = 12'h00f;
rom[788] = 12'h000;
rom[789] = 12'h000;
rom[790] = 12'h000;
rom[791] = 12'h000;
rom[792] = 12'h000;
rom[793] = 12'h000;
rom[794] = 12'h000;
rom[795] = 12'h000;
rom[796] = 12'h000;
rom[797] = 12'h000;
rom[798] = 12'h000;
rom[799] = 12'h000;
rom[800] = 12'h007;
rom[801] = 12'h007;
rom[802] = 12'h000;
rom[803] = 12'h000;
rom[804] = 12'h000;
rom[805] = 12'h000;
rom[806] = 12'h000;
rom[807] = 12'h000;
rom[808] = 12'h00f;
rom[809] = 12'h00f;
rom[810] = 12'h00f;
rom[811] = 12'h00f;
rom[812] = 12'h00f;
rom[813] = 12'h00f;
rom[814] = 12'h000;
rom[815] = 12'h000;
rom[816] = 12'h000;
rom[817] = 12'h000;
rom[818] = 12'h000;
rom[819] = 12'h000;
rom[820] = 12'h000;
rom[821] = 12'h000;
rom[822] = 12'h000;
rom[823] = 12'h000;
rom[824] = 12'h000;
rom[825] = 12'h000;
rom[826] = 12'h007;
rom[827] = 12'h007;
rom[828] = 12'h000;
rom[829] = 12'h000;
rom[830] = 12'h000;
rom[831] = 12'h000;
rom[832] = 12'h000;
rom[833] = 12'h000;
rom[834] = 12'h00f;
rom[835] = 12'h00f;
rom[836] = 12'h00f;
rom[837] = 12'h00f;
rom[838] = 12'h00f;
rom[839] = 12'h00f;
rom[840] = 12'h000;
rom[841] = 12'h000;
rom[842] = 12'h000;
rom[843] = 12'h000;
rom[844] = 12'h000;
rom[845] = 12'h000;
rom[846] = 12'h000;
rom[847] = 12'h000;
rom[848] = 12'h000;
rom[849] = 12'h000;
rom[850] = 12'h007;
rom[851] = 12'h007;
rom[852] = 12'h000;
rom[853] = 12'h000;
rom[854] = 12'h007;
rom[855] = 12'h007;
rom[856] = 12'h000;
rom[857] = 12'h000;
rom[858] = 12'h000;
rom[859] = 12'h000;
rom[860] = 12'h00f;
rom[861] = 12'h00f;
rom[862] = 12'h00f;
rom[863] = 12'h00f;
rom[864] = 12'h00f;
rom[865] = 12'h00f;
rom[866] = 12'h000;
rom[867] = 12'h000;
rom[868] = 12'h000;
rom[869] = 12'h000;
rom[870] = 12'h000;
rom[871] = 12'h000;
rom[872] = 12'h000;
rom[873] = 12'h000;
rom[874] = 12'h000;
rom[875] = 12'h000;
rom[876] = 12'h007;
rom[877] = 12'h007;
rom[878] = 12'h000;
rom[879] = 12'h000;
rom[880] = 12'h007;
rom[881] = 12'h007;
rom[882] = 12'h000;
rom[883] = 12'h000;
rom[884] = 12'h000;
rom[885] = 12'h000;
rom[886] = 12'h00f;
rom[887] = 12'h00f;
rom[888] = 12'h00f;
rom[889] = 12'h00f;
rom[890] = 12'h00f;
rom[891] = 12'h00f;
rom[892] = 12'h000;
rom[893] = 12'h000;
rom[894] = 12'h000;
rom[895] = 12'h000;
rom[896] = 12'h000;
rom[897] = 12'h000;
rom[898] = 12'h000;
rom[899] = 12'h000;
rom[900] = 12'h000;
rom[901] = 12'h000;
rom[902] = 12'h000;
rom[903] = 12'h000;
rom[904] = 12'h007;
rom[905] = 12'h007;
rom[906] = 12'h000;
rom[907] = 12'h000;
rom[908] = 12'h000;
rom[909] = 12'h000;
rom[910] = 12'h000;
rom[911] = 12'h000;
rom[912] = 12'h00f;
rom[913] = 12'h00f;
rom[914] = 12'h00f;
rom[915] = 12'h00f;
rom[916] = 12'h00f;
rom[917] = 12'h00f;
rom[918] = 12'h000;
rom[919] = 12'h000;
rom[920] = 12'h000;
rom[921] = 12'h000;
rom[922] = 12'h000;
rom[923] = 12'h000;
rom[924] = 12'h000;
rom[925] = 12'h000;
rom[926] = 12'h000;
rom[927] = 12'h000;
rom[928] = 12'h000;
rom[929] = 12'h000;
rom[930] = 12'h007;
rom[931] = 12'h007;
rom[932] = 12'h000;
rom[933] = 12'h000;
rom[934] = 12'h000;
rom[935] = 12'h000;
rom[936] = 12'h000;
rom[937] = 12'h000;
rom[938] = 12'h00f;
rom[939] = 12'h00f;
rom[940] = 12'h00f;
rom[941] = 12'h00f;
rom[942] = 12'h00f;
rom[943] = 12'h00f;
rom[944] = 12'h000;
rom[945] = 12'h000;
rom[946] = 12'h000;
rom[947] = 12'h000;
rom[948] = 12'h000;
rom[949] = 12'h000;
rom[950] = 12'h000;
rom[951] = 12'h000;
rom[952] = 12'h000;
rom[953] = 12'h000;
rom[954] = 12'h007;
rom[955] = 12'h007;
rom[956] = 12'h000;
rom[957] = 12'h000;
rom[958] = 12'h007;
rom[959] = 12'h007;
rom[960] = 12'h000;
rom[961] = 12'h000;
rom[962] = 12'h000;
rom[963] = 12'h000;
rom[964] = 12'h00f;
rom[965] = 12'h00f;
rom[966] = 12'h00f;
rom[967] = 12'h00f;
rom[968] = 12'h00f;
rom[969] = 12'h00f;
rom[970] = 12'h000;
rom[971] = 12'h000;
rom[972] = 12'h000;
rom[973] = 12'h000;
rom[974] = 12'h000;
rom[975] = 12'h000;
rom[976] = 12'h000;
rom[977] = 12'h000;
rom[978] = 12'h000;
rom[979] = 12'h000;
rom[980] = 12'h007;
rom[981] = 12'h007;
rom[982] = 12'h000;
rom[983] = 12'h000;
rom[984] = 12'h007;
rom[985] = 12'h007;
rom[986] = 12'h000;
rom[987] = 12'h000;
rom[988] = 12'h000;
rom[989] = 12'h000;
rom[990] = 12'h00f;
rom[991] = 12'h00f;
rom[992] = 12'h00f;
rom[993] = 12'h00f;
rom[994] = 12'h000;
rom[995] = 12'h000;
rom[996] = 12'h00f;
rom[997] = 12'h00f;
rom[998] = 12'h00f;
rom[999] = 12'h00f;
rom[1000] = 12'h00f;
rom[1001] = 12'h00f;
rom[1002] = 12'h00f;
rom[1003] = 12'h00f;
rom[1004] = 12'h00f;
rom[1005] = 12'h00f;
rom[1006] = 12'h000;
rom[1007] = 12'h000;
rom[1008] = 12'h007;
rom[1009] = 12'h007;
rom[1010] = 12'h000;
rom[1011] = 12'h000;
rom[1012] = 12'h000;
rom[1013] = 12'h000;
rom[1014] = 12'h000;
rom[1015] = 12'h000;
rom[1016] = 12'h00f;
rom[1017] = 12'h00f;
rom[1018] = 12'h00f;
rom[1019] = 12'h00f;
rom[1020] = 12'h000;
rom[1021] = 12'h000;
rom[1022] = 12'h00f;
rom[1023] = 12'h00f;
rom[1024] = 12'h00f;
rom[1025] = 12'h00f;
rom[1026] = 12'h00f;
rom[1027] = 12'h00f;
rom[1028] = 12'h00f;
rom[1029] = 12'h00f;
rom[1030] = 12'h00f;
rom[1031] = 12'h00f;
rom[1032] = 12'h000;
rom[1033] = 12'h000;
rom[1034] = 12'h007;
rom[1035] = 12'h007;
rom[1036] = 12'h000;
rom[1037] = 12'h000;
rom[1038] = 12'h000;
rom[1039] = 12'h000;
rom[1040] = 12'h000;
rom[1041] = 12'h000;
rom[1042] = 12'h00f;
rom[1043] = 12'h00f;
rom[1044] = 12'h000;
rom[1045] = 12'h000;
rom[1046] = 12'h00f;
rom[1047] = 12'h00f;
rom[1048] = 12'h00f;
rom[1049] = 12'h00f;
rom[1050] = 12'h00f;
rom[1051] = 12'h00f;
rom[1052] = 12'h00f;
rom[1053] = 12'h00f;
rom[1054] = 12'h00f;
rom[1055] = 12'h00f;
rom[1056] = 12'h00f;
rom[1057] = 12'h00f;
rom[1058] = 12'h00f;
rom[1059] = 12'h00f;
rom[1060] = 12'h000;
rom[1061] = 12'h000;
rom[1062] = 12'h007;
rom[1063] = 12'h007;
rom[1064] = 12'h000;
rom[1065] = 12'h000;
rom[1066] = 12'h000;
rom[1067] = 12'h000;
rom[1068] = 12'h00f;
rom[1069] = 12'h00f;
rom[1070] = 12'h000;
rom[1071] = 12'h000;
rom[1072] = 12'h00f;
rom[1073] = 12'h00f;
rom[1074] = 12'h00f;
rom[1075] = 12'h00f;
rom[1076] = 12'h00f;
rom[1077] = 12'h00f;
rom[1078] = 12'h00f;
rom[1079] = 12'h00f;
rom[1080] = 12'h00f;
rom[1081] = 12'h00f;
rom[1082] = 12'h00f;
rom[1083] = 12'h00f;
rom[1084] = 12'h00f;
rom[1085] = 12'h00f;
rom[1086] = 12'h000;
rom[1087] = 12'h000;
rom[1088] = 12'h007;
rom[1089] = 12'h007;
rom[1090] = 12'h000;
rom[1091] = 12'h000;
rom[1092] = 12'h000;
rom[1093] = 12'h000;
rom[1094] = 12'h000;
rom[1095] = 12'h000;
rom[1096] = 12'h00f;
rom[1097] = 12'h00f;
rom[1098] = 12'h00f;
rom[1099] = 12'h00f;
rom[1100] = 12'h00f;
rom[1101] = 12'h00f;
rom[1102] = 12'h00f;
rom[1103] = 12'h00f;
rom[1104] = 12'h00f;
rom[1105] = 12'h00f;
rom[1106] = 12'h00f;
rom[1107] = 12'h00f;
rom[1108] = 12'h00f;
rom[1109] = 12'h00f;
rom[1110] = 12'h00f;
rom[1111] = 12'h00f;
rom[1112] = 12'h00f;
rom[1113] = 12'h00f;
rom[1114] = 12'h000;
rom[1115] = 12'h000;
rom[1116] = 12'h000;
rom[1117] = 12'h000;
rom[1118] = 12'h000;
rom[1119] = 12'h000;
rom[1120] = 12'h000;
rom[1121] = 12'h000;
rom[1122] = 12'h00f;
rom[1123] = 12'h00f;
rom[1124] = 12'h00f;
rom[1125] = 12'h00f;
rom[1126] = 12'h00f;
rom[1127] = 12'h00f;
rom[1128] = 12'h00f;
rom[1129] = 12'h00f;
rom[1130] = 12'h00f;
rom[1131] = 12'h00f;
rom[1132] = 12'h00f;
rom[1133] = 12'h00f;
rom[1134] = 12'h00f;
rom[1135] = 12'h00f;
rom[1136] = 12'h00f;
rom[1137] = 12'h00f;
rom[1138] = 12'h00f;
rom[1139] = 12'h00f;
rom[1140] = 12'h000;
rom[1141] = 12'h000;
rom[1142] = 12'h000;
rom[1143] = 12'h000;
rom[1144] = 12'h000;
rom[1145] = 12'h000;
rom[1146] = 12'h000;
rom[1147] = 12'h000;
rom[1148] = 12'h000;
rom[1149] = 12'h000;
rom[1150] = 12'h000;
rom[1151] = 12'h000;
rom[1152] = 12'h000;
rom[1153] = 12'h000;
rom[1154] = 12'h000;
rom[1155] = 12'h000;
rom[1156] = 12'h000;
rom[1157] = 12'h000;
rom[1158] = 12'h000;
rom[1159] = 12'h000;
rom[1160] = 12'h000;
rom[1161] = 12'h000;
rom[1162] = 12'h000;
rom[1163] = 12'h000;
rom[1164] = 12'h000;
rom[1165] = 12'h000;
rom[1166] = 12'h000;
rom[1167] = 12'h000;
rom[1168] = 12'h000;
rom[1169] = 12'h000;
rom[1170] = 12'h000;
rom[1171] = 12'h000;
rom[1172] = 12'h000;
rom[1173] = 12'h000;
rom[1174] = 12'h000;
rom[1175] = 12'h000;
rom[1176] = 12'h000;
rom[1177] = 12'h000;
rom[1178] = 12'h000;
rom[1179] = 12'h000;
rom[1180] = 12'h000;
rom[1181] = 12'h000;
rom[1182] = 12'h000;
rom[1183] = 12'h000;
rom[1184] = 12'h000;
rom[1185] = 12'h000;
rom[1186] = 12'h000;
rom[1187] = 12'h000;
rom[1188] = 12'h000;
rom[1189] = 12'h000;
rom[1190] = 12'h000;
rom[1191] = 12'h000;
rom[1192] = 12'h000;
rom[1193] = 12'h000;
rom[1194] = 12'h000;
rom[1195] = 12'h000;
  end
  endmodule

    module dash_rom (                       //три
  input  wire    [13:0]     addr,
  output wire    [11:0]     word
);

  logic [11:0] rom [(46 * 26)];

  assign word = rom[addr];

  initial begin
rom[0] = 12'h000;
rom[1] = 12'h000;
rom[2] = 12'h000;
rom[3] = 12'h000;
rom[4] = 12'h000;
rom[5] = 12'h000;
rom[6] = 12'h000;
rom[7] = 12'h000;
rom[8] = 12'h000;
rom[9] = 12'h000;
rom[10] = 12'h000;
rom[11] = 12'h000;
rom[12] = 12'h000;
rom[13] = 12'h000;
rom[14] = 12'h000;
rom[15] = 12'h000;
rom[16] = 12'h000;
rom[17] = 12'h000;
rom[18] = 12'h000;
rom[19] = 12'h000;
rom[20] = 12'h000;
rom[21] = 12'h000;
rom[22] = 12'h000;
rom[23] = 12'h000;
rom[24] = 12'h000;
rom[25] = 12'h000;
rom[26] = 12'h000;
rom[27] = 12'h000;
rom[28] = 12'h000;
rom[29] = 12'h000;
rom[30] = 12'h000;
rom[31] = 12'h000;
rom[32] = 12'h000;
rom[33] = 12'h000;
rom[34] = 12'h000;
rom[35] = 12'h000;
rom[36] = 12'h000;
rom[37] = 12'h000;
rom[38] = 12'h000;
rom[39] = 12'h000;
rom[40] = 12'h000;
rom[41] = 12'h000;
rom[42] = 12'h000;
rom[43] = 12'h000;
rom[44] = 12'h000;
rom[45] = 12'h000;
rom[46] = 12'h000;
rom[47] = 12'h000;
rom[48] = 12'h000;
rom[49] = 12'h000;
rom[50] = 12'h000;
rom[51] = 12'h000;
rom[52] = 12'h000;
rom[53] = 12'h000;
rom[54] = 12'h000;
rom[55] = 12'h000;
rom[56] = 12'h00f;
rom[57] = 12'h00f;
rom[58] = 12'h00f;
rom[59] = 12'h00f;
rom[60] = 12'h00f;
rom[61] = 12'h00f;
rom[62] = 12'h00f;
rom[63] = 12'h00f;
rom[64] = 12'h00f;
rom[65] = 12'h00f;
rom[66] = 12'h00f;
rom[67] = 12'h00f;
rom[68] = 12'h00f;
rom[69] = 12'h00f;
rom[70] = 12'h00f;
rom[71] = 12'h00f;
rom[72] = 12'h00f;
rom[73] = 12'h00f;
rom[74] = 12'h000;
rom[75] = 12'h000;
rom[76] = 12'h000;
rom[77] = 12'h000;
rom[78] = 12'h000;
rom[79] = 12'h000;
rom[80] = 12'h000;
rom[81] = 12'h000;
rom[82] = 12'h00f;
rom[83] = 12'h00f;
rom[84] = 12'h00f;
rom[85] = 12'h00f;
rom[86] = 12'h00f;
rom[87] = 12'h00f;
rom[88] = 12'h00f;
rom[89] = 12'h00f;
rom[90] = 12'h00f;
rom[91] = 12'h00f;
rom[92] = 12'h00f;
rom[93] = 12'h00f;
rom[94] = 12'h00f;
rom[95] = 12'h00f;
rom[96] = 12'h00f;
rom[97] = 12'h00f;
rom[98] = 12'h00f;
rom[99] = 12'h00f;
rom[100] = 12'h000;
rom[101] = 12'h000;
rom[102] = 12'h000;
rom[103] = 12'h000;
rom[104] = 12'h000;
rom[105] = 12'h000;
rom[106] = 12'h007;
rom[107] = 12'h007;
rom[108] = 12'h000;
rom[109] = 12'h000;
rom[110] = 12'h00f;
rom[111] = 12'h00f;
rom[112] = 12'h00f;
rom[113] = 12'h00f;
rom[114] = 12'h00f;
rom[115] = 12'h00f;
rom[116] = 12'h00f;
rom[117] = 12'h00f;
rom[118] = 12'h00f;
rom[119] = 12'h00f;
rom[120] = 12'h00f;
rom[121] = 12'h00f;
rom[122] = 12'h00f;
rom[123] = 12'h00f;
rom[124] = 12'h000;
rom[125] = 12'h000;
rom[126] = 12'h00f;
rom[127] = 12'h00f;
rom[128] = 12'h000;
rom[129] = 12'h000;
rom[130] = 12'h000;
rom[131] = 12'h000;
rom[132] = 12'h007;
rom[133] = 12'h007;
rom[134] = 12'h000;
rom[135] = 12'h000;
rom[136] = 12'h00f;
rom[137] = 12'h00f;
rom[138] = 12'h00f;
rom[139] = 12'h00f;
rom[140] = 12'h00f;
rom[141] = 12'h00f;
rom[142] = 12'h00f;
rom[143] = 12'h00f;
rom[144] = 12'h00f;
rom[145] = 12'h00f;
rom[146] = 12'h00f;
rom[147] = 12'h00f;
rom[148] = 12'h00f;
rom[149] = 12'h00f;
rom[150] = 12'h000;
rom[151] = 12'h000;
rom[152] = 12'h00f;
rom[153] = 12'h00f;
rom[154] = 12'h000;
rom[155] = 12'h000;
rom[156] = 12'h000;
rom[157] = 12'h000;
rom[158] = 12'h000;
rom[159] = 12'h000;
rom[160] = 12'h007;
rom[161] = 12'h007;
rom[162] = 12'h000;
rom[163] = 12'h000;
rom[164] = 12'h00f;
rom[165] = 12'h00f;
rom[166] = 12'h00f;
rom[167] = 12'h00f;
rom[168] = 12'h00f;
rom[169] = 12'h00f;
rom[170] = 12'h00f;
rom[171] = 12'h00f;
rom[172] = 12'h00f;
rom[173] = 12'h00f;
rom[174] = 12'h000;
rom[175] = 12'h000;
rom[176] = 12'h00f;
rom[177] = 12'h00f;
rom[178] = 12'h00f;
rom[179] = 12'h00f;
rom[180] = 12'h000;
rom[181] = 12'h000;
rom[182] = 12'h000;
rom[183] = 12'h000;
rom[184] = 12'h000;
rom[185] = 12'h000;
rom[186] = 12'h007;
rom[187] = 12'h007;
rom[188] = 12'h000;
rom[189] = 12'h000;
rom[190] = 12'h00f;
rom[191] = 12'h00f;
rom[192] = 12'h00f;
rom[193] = 12'h00f;
rom[194] = 12'h00f;
rom[195] = 12'h00f;
rom[196] = 12'h00f;
rom[197] = 12'h00f;
rom[198] = 12'h00f;
rom[199] = 12'h00f;
rom[200] = 12'h000;
rom[201] = 12'h000;
rom[202] = 12'h00f;
rom[203] = 12'h00f;
rom[204] = 12'h00f;
rom[205] = 12'h00f;
rom[206] = 12'h000;
rom[207] = 12'h000;
rom[208] = 12'h000;
rom[209] = 12'h000;
rom[210] = 12'h007;
rom[211] = 12'h007;
rom[212] = 12'h000;
rom[213] = 12'h000;
rom[214] = 12'h007;
rom[215] = 12'h007;
rom[216] = 12'h000;
rom[217] = 12'h000;
rom[218] = 12'h000;
rom[219] = 12'h000;
rom[220] = 12'h000;
rom[221] = 12'h000;
rom[222] = 12'h000;
rom[223] = 12'h000;
rom[224] = 12'h000;
rom[225] = 12'h000;
rom[226] = 12'h00f;
rom[227] = 12'h00f;
rom[228] = 12'h00f;
rom[229] = 12'h00f;
rom[230] = 12'h00f;
rom[231] = 12'h00f;
rom[232] = 12'h000;
rom[233] = 12'h000;
rom[234] = 12'h000;
rom[235] = 12'h000;
rom[236] = 12'h007;
rom[237] = 12'h007;
rom[238] = 12'h000;
rom[239] = 12'h000;
rom[240] = 12'h007;
rom[241] = 12'h007;
rom[242] = 12'h000;
rom[243] = 12'h000;
rom[244] = 12'h000;
rom[245] = 12'h000;
rom[246] = 12'h000;
rom[247] = 12'h000;
rom[248] = 12'h000;
rom[249] = 12'h000;
rom[250] = 12'h000;
rom[251] = 12'h000;
rom[252] = 12'h00f;
rom[253] = 12'h00f;
rom[254] = 12'h00f;
rom[255] = 12'h00f;
rom[256] = 12'h00f;
rom[257] = 12'h00f;
rom[258] = 12'h000;
rom[259] = 12'h000;
rom[260] = 12'h000;
rom[261] = 12'h000;
rom[262] = 12'h000;
rom[263] = 12'h000;
rom[264] = 12'h007;
rom[265] = 12'h007;
rom[266] = 12'h000;
rom[267] = 12'h000;
rom[268] = 12'h000;
rom[269] = 12'h000;
rom[270] = 12'h000;
rom[271] = 12'h000;
rom[272] = 12'h000;
rom[273] = 12'h000;
rom[274] = 12'h000;
rom[275] = 12'h000;
rom[276] = 12'h000;
rom[277] = 12'h000;
rom[278] = 12'h00f;
rom[279] = 12'h00f;
rom[280] = 12'h00f;
rom[281] = 12'h00f;
rom[282] = 12'h00f;
rom[283] = 12'h00f;
rom[284] = 12'h000;
rom[285] = 12'h000;
rom[286] = 12'h000;
rom[287] = 12'h000;
rom[288] = 12'h000;
rom[289] = 12'h000;
rom[290] = 12'h007;
rom[291] = 12'h007;
rom[292] = 12'h000;
rom[293] = 12'h000;
rom[294] = 12'h000;
rom[295] = 12'h000;
rom[296] = 12'h000;
rom[297] = 12'h000;
rom[298] = 12'h000;
rom[299] = 12'h000;
rom[300] = 12'h000;
rom[301] = 12'h000;
rom[302] = 12'h000;
rom[303] = 12'h000;
rom[304] = 12'h00f;
rom[305] = 12'h00f;
rom[306] = 12'h00f;
rom[307] = 12'h00f;
rom[308] = 12'h00f;
rom[309] = 12'h00f;
rom[310] = 12'h000;
rom[311] = 12'h000;
rom[312] = 12'h000;
rom[313] = 12'h000;
rom[314] = 12'h007;
rom[315] = 12'h007;
rom[316] = 12'h000;
rom[317] = 12'h000;
rom[318] = 12'h007;
rom[319] = 12'h007;
rom[320] = 12'h000;
rom[321] = 12'h000;
rom[322] = 12'h000;
rom[323] = 12'h000;
rom[324] = 12'h000;
rom[325] = 12'h000;
rom[326] = 12'h000;
rom[327] = 12'h000;
rom[328] = 12'h000;
rom[329] = 12'h000;
rom[330] = 12'h00f;
rom[331] = 12'h00f;
rom[332] = 12'h00f;
rom[333] = 12'h00f;
rom[334] = 12'h00f;
rom[335] = 12'h00f;
rom[336] = 12'h000;
rom[337] = 12'h000;
rom[338] = 12'h000;
rom[339] = 12'h000;
rom[340] = 12'h007;
rom[341] = 12'h007;
rom[342] = 12'h000;
rom[343] = 12'h000;
rom[344] = 12'h007;
rom[345] = 12'h007;
rom[346] = 12'h000;
rom[347] = 12'h000;
rom[348] = 12'h000;
rom[349] = 12'h000;
rom[350] = 12'h000;
rom[351] = 12'h000;
rom[352] = 12'h000;
rom[353] = 12'h000;
rom[354] = 12'h000;
rom[355] = 12'h000;
rom[356] = 12'h00f;
rom[357] = 12'h00f;
rom[358] = 12'h00f;
rom[359] = 12'h00f;
rom[360] = 12'h00f;
rom[361] = 12'h00f;
rom[362] = 12'h000;
rom[363] = 12'h000;
rom[364] = 12'h000;
rom[365] = 12'h000;
rom[366] = 12'h000;
rom[367] = 12'h000;
rom[368] = 12'h007;
rom[369] = 12'h007;
rom[370] = 12'h000;
rom[371] = 12'h000;
rom[372] = 12'h000;
rom[373] = 12'h000;
rom[374] = 12'h000;
rom[375] = 12'h000;
rom[376] = 12'h000;
rom[377] = 12'h000;
rom[378] = 12'h000;
rom[379] = 12'h000;
rom[380] = 12'h000;
rom[381] = 12'h000;
rom[382] = 12'h00f;
rom[383] = 12'h00f;
rom[384] = 12'h00f;
rom[385] = 12'h00f;
rom[386] = 12'h00f;
rom[387] = 12'h00f;
rom[388] = 12'h000;
rom[389] = 12'h000;
rom[390] = 12'h000;
rom[391] = 12'h000;
rom[392] = 12'h000;
rom[393] = 12'h000;
rom[394] = 12'h007;
rom[395] = 12'h007;
rom[396] = 12'h000;
rom[397] = 12'h000;
rom[398] = 12'h000;
rom[399] = 12'h000;
rom[400] = 12'h000;
rom[401] = 12'h000;
rom[402] = 12'h000;
rom[403] = 12'h000;
rom[404] = 12'h000;
rom[405] = 12'h000;
rom[406] = 12'h000;
rom[407] = 12'h000;
rom[408] = 12'h00f;
rom[409] = 12'h00f;
rom[410] = 12'h00f;
rom[411] = 12'h00f;
rom[412] = 12'h00f;
rom[413] = 12'h00f;
rom[414] = 12'h000;
rom[415] = 12'h000;
rom[416] = 12'h000;
rom[417] = 12'h000;
rom[418] = 12'h007;
rom[419] = 12'h007;
rom[420] = 12'h000;
rom[421] = 12'h000;
rom[422] = 12'h007;
rom[423] = 12'h007;
rom[424] = 12'h000;
rom[425] = 12'h000;
rom[426] = 12'h000;
rom[427] = 12'h000;
rom[428] = 12'h000;
rom[429] = 12'h000;
rom[430] = 12'h000;
rom[431] = 12'h000;
rom[432] = 12'h000;
rom[433] = 12'h000;
rom[434] = 12'h00f;
rom[435] = 12'h00f;
rom[436] = 12'h00f;
rom[437] = 12'h00f;
rom[438] = 12'h00f;
rom[439] = 12'h00f;
rom[440] = 12'h000;
rom[441] = 12'h000;
rom[442] = 12'h000;
rom[443] = 12'h000;
rom[444] = 12'h007;
rom[445] = 12'h007;
rom[446] = 12'h000;
rom[447] = 12'h000;
rom[448] = 12'h007;
rom[449] = 12'h007;
rom[450] = 12'h000;
rom[451] = 12'h000;
rom[452] = 12'h000;
rom[453] = 12'h000;
rom[454] = 12'h000;
rom[455] = 12'h000;
rom[456] = 12'h000;
rom[457] = 12'h000;
rom[458] = 12'h000;
rom[459] = 12'h000;
rom[460] = 12'h00f;
rom[461] = 12'h00f;
rom[462] = 12'h00f;
rom[463] = 12'h00f;
rom[464] = 12'h00f;
rom[465] = 12'h00f;
rom[466] = 12'h000;
rom[467] = 12'h000;
rom[468] = 12'h000;
rom[469] = 12'h000;
rom[470] = 12'h000;
rom[471] = 12'h000;
rom[472] = 12'h007;
rom[473] = 12'h007;
rom[474] = 12'h000;
rom[475] = 12'h000;
rom[476] = 12'h000;
rom[477] = 12'h000;
rom[478] = 12'h000;
rom[479] = 12'h000;
rom[480] = 12'h000;
rom[481] = 12'h000;
rom[482] = 12'h000;
rom[483] = 12'h000;
rom[484] = 12'h000;
rom[485] = 12'h000;
rom[486] = 12'h000;
rom[487] = 12'h000;
rom[488] = 12'h00f;
rom[489] = 12'h00f;
rom[490] = 12'h00f;
rom[491] = 12'h00f;
rom[492] = 12'h000;
rom[493] = 12'h000;
rom[494] = 12'h000;
rom[495] = 12'h000;
rom[496] = 12'h000;
rom[497] = 12'h000;
rom[498] = 12'h007;
rom[499] = 12'h007;
rom[500] = 12'h000;
rom[501] = 12'h000;
rom[502] = 12'h000;
rom[503] = 12'h000;
rom[504] = 12'h000;
rom[505] = 12'h000;
rom[506] = 12'h000;
rom[507] = 12'h000;
rom[508] = 12'h000;
rom[509] = 12'h000;
rom[510] = 12'h000;
rom[511] = 12'h000;
rom[512] = 12'h000;
rom[513] = 12'h000;
rom[514] = 12'h00f;
rom[515] = 12'h00f;
rom[516] = 12'h00f;
rom[517] = 12'h00f;
rom[518] = 12'h000;
rom[519] = 12'h000;
rom[520] = 12'h000;
rom[521] = 12'h000;
rom[522] = 12'h007;
rom[523] = 12'h007;
rom[524] = 12'h000;
rom[525] = 12'h000;
rom[526] = 12'h00f;
rom[527] = 12'h00f;
rom[528] = 12'h00f;
rom[529] = 12'h00f;
rom[530] = 12'h00f;
rom[531] = 12'h00f;
rom[532] = 12'h00f;
rom[533] = 12'h00f;
rom[534] = 12'h00f;
rom[535] = 12'h00f;
rom[536] = 12'h00f;
rom[537] = 12'h00f;
rom[538] = 12'h00f;
rom[539] = 12'h00f;
rom[540] = 12'h000;
rom[541] = 12'h000;
rom[542] = 12'h00f;
rom[543] = 12'h00f;
rom[544] = 12'h000;
rom[545] = 12'h000;
rom[546] = 12'h000;
rom[547] = 12'h000;
rom[548] = 12'h007;
rom[549] = 12'h007;
rom[550] = 12'h000;
rom[551] = 12'h000;
rom[552] = 12'h00f;
rom[553] = 12'h00f;
rom[554] = 12'h00f;
rom[555] = 12'h00f;
rom[556] = 12'h00f;
rom[557] = 12'h00f;
rom[558] = 12'h00f;
rom[559] = 12'h00f;
rom[560] = 12'h00f;
rom[561] = 12'h00f;
rom[562] = 12'h00f;
rom[563] = 12'h00f;
rom[564] = 12'h00f;
rom[565] = 12'h00f;
rom[566] = 12'h000;
rom[567] = 12'h000;
rom[568] = 12'h00f;
rom[569] = 12'h00f;
rom[570] = 12'h000;
rom[571] = 12'h000;
rom[572] = 12'h000;
rom[573] = 12'h000;
rom[574] = 12'h000;
rom[575] = 12'h000;
rom[576] = 12'h00f;
rom[577] = 12'h00f;
rom[578] = 12'h00f;
rom[579] = 12'h00f;
rom[580] = 12'h00f;
rom[581] = 12'h00f;
rom[582] = 12'h00f;
rom[583] = 12'h00f;
rom[584] = 12'h00f;
rom[585] = 12'h00f;
rom[586] = 12'h00f;
rom[587] = 12'h00f;
rom[588] = 12'h00f;
rom[589] = 12'h00f;
rom[590] = 12'h00f;
rom[591] = 12'h00f;
rom[592] = 12'h00f;
rom[593] = 12'h00f;
rom[594] = 12'h000;
rom[595] = 12'h000;
rom[596] = 12'h000;
rom[597] = 12'h000;
rom[598] = 12'h000;
rom[599] = 12'h000;
rom[600] = 12'h000;
rom[601] = 12'h000;
rom[602] = 12'h00f;
rom[603] = 12'h00f;
rom[604] = 12'h00f;
rom[605] = 12'h00f;
rom[606] = 12'h00f;
rom[607] = 12'h00f;
rom[608] = 12'h00f;
rom[609] = 12'h00f;
rom[610] = 12'h00f;
rom[611] = 12'h00f;
rom[612] = 12'h00f;
rom[613] = 12'h00f;
rom[614] = 12'h00f;
rom[615] = 12'h00f;
rom[616] = 12'h00f;
rom[617] = 12'h00f;
rom[618] = 12'h00f;
rom[619] = 12'h00f;
rom[620] = 12'h000;
rom[621] = 12'h000;
rom[622] = 12'h000;
rom[623] = 12'h000;
rom[624] = 12'h000;
rom[625] = 12'h000;
rom[626] = 12'h007;
rom[627] = 12'h007;
rom[628] = 12'h000;
rom[629] = 12'h000;
rom[630] = 12'h00f;
rom[631] = 12'h00f;
rom[632] = 12'h00f;
rom[633] = 12'h00f;
rom[634] = 12'h00f;
rom[635] = 12'h00f;
rom[636] = 12'h00f;
rom[637] = 12'h00f;
rom[638] = 12'h00f;
rom[639] = 12'h00f;
rom[640] = 12'h00f;
rom[641] = 12'h00f;
rom[642] = 12'h00f;
rom[643] = 12'h00f;
rom[644] = 12'h000;
rom[645] = 12'h000;
rom[646] = 12'h00f;
rom[647] = 12'h00f;
rom[648] = 12'h000;
rom[649] = 12'h000;
rom[650] = 12'h000;
rom[651] = 12'h000;
rom[652] = 12'h007;
rom[653] = 12'h007;
rom[654] = 12'h000;
rom[655] = 12'h000;
rom[656] = 12'h00f;
rom[657] = 12'h00f;
rom[658] = 12'h00f;
rom[659] = 12'h00f;
rom[660] = 12'h00f;
rom[661] = 12'h00f;
rom[662] = 12'h00f;
rom[663] = 12'h00f;
rom[664] = 12'h00f;
rom[665] = 12'h00f;
rom[666] = 12'h00f;
rom[667] = 12'h00f;
rom[668] = 12'h00f;
rom[669] = 12'h00f;
rom[670] = 12'h000;
rom[671] = 12'h000;
rom[672] = 12'h00f;
rom[673] = 12'h00f;
rom[674] = 12'h000;
rom[675] = 12'h000;
rom[676] = 12'h000;
rom[677] = 12'h000;
rom[678] = 12'h000;
rom[679] = 12'h000;
rom[680] = 12'h007;
rom[681] = 12'h007;
rom[682] = 12'h000;
rom[683] = 12'h000;
rom[684] = 12'h000;
rom[685] = 12'h000;
rom[686] = 12'h000;
rom[687] = 12'h000;
rom[688] = 12'h000;
rom[689] = 12'h000;
rom[690] = 12'h000;
rom[691] = 12'h000;
rom[692] = 12'h000;
rom[693] = 12'h000;
rom[694] = 12'h000;
rom[695] = 12'h000;
rom[696] = 12'h00f;
rom[697] = 12'h00f;
rom[698] = 12'h00f;
rom[699] = 12'h00f;
rom[700] = 12'h000;
rom[701] = 12'h000;
rom[702] = 12'h000;
rom[703] = 12'h000;
rom[704] = 12'h000;
rom[705] = 12'h000;
rom[706] = 12'h007;
rom[707] = 12'h007;
rom[708] = 12'h000;
rom[709] = 12'h000;
rom[710] = 12'h000;
rom[711] = 12'h000;
rom[712] = 12'h000;
rom[713] = 12'h000;
rom[714] = 12'h000;
rom[715] = 12'h000;
rom[716] = 12'h000;
rom[717] = 12'h000;
rom[718] = 12'h000;
rom[719] = 12'h000;
rom[720] = 12'h000;
rom[721] = 12'h000;
rom[722] = 12'h00f;
rom[723] = 12'h00f;
rom[724] = 12'h00f;
rom[725] = 12'h00f;
rom[726] = 12'h000;
rom[727] = 12'h000;
rom[728] = 12'h000;
rom[729] = 12'h000;
rom[730] = 12'h007;
rom[731] = 12'h007;
rom[732] = 12'h000;
rom[733] = 12'h000;
rom[734] = 12'h007;
rom[735] = 12'h007;
rom[736] = 12'h000;
rom[737] = 12'h000;
rom[738] = 12'h000;
rom[739] = 12'h000;
rom[740] = 12'h000;
rom[741] = 12'h000;
rom[742] = 12'h000;
rom[743] = 12'h000;
rom[744] = 12'h000;
rom[745] = 12'h000;
rom[746] = 12'h00f;
rom[747] = 12'h00f;
rom[748] = 12'h00f;
rom[749] = 12'h00f;
rom[750] = 12'h00f;
rom[751] = 12'h00f;
rom[752] = 12'h000;
rom[753] = 12'h000;
rom[754] = 12'h000;
rom[755] = 12'h000;
rom[756] = 12'h007;
rom[757] = 12'h007;
rom[758] = 12'h000;
rom[759] = 12'h000;
rom[760] = 12'h007;
rom[761] = 12'h007;
rom[762] = 12'h000;
rom[763] = 12'h000;
rom[764] = 12'h000;
rom[765] = 12'h000;
rom[766] = 12'h000;
rom[767] = 12'h000;
rom[768] = 12'h000;
rom[769] = 12'h000;
rom[770] = 12'h000;
rom[771] = 12'h000;
rom[772] = 12'h00f;
rom[773] = 12'h00f;
rom[774] = 12'h00f;
rom[775] = 12'h00f;
rom[776] = 12'h00f;
rom[777] = 12'h00f;
rom[778] = 12'h000;
rom[779] = 12'h000;
rom[780] = 12'h000;
rom[781] = 12'h000;
rom[782] = 12'h000;
rom[783] = 12'h000;
rom[784] = 12'h007;
rom[785] = 12'h007;
rom[786] = 12'h000;
rom[787] = 12'h000;
rom[788] = 12'h000;
rom[789] = 12'h000;
rom[790] = 12'h000;
rom[791] = 12'h000;
rom[792] = 12'h000;
rom[793] = 12'h000;
rom[794] = 12'h000;
rom[795] = 12'h000;
rom[796] = 12'h000;
rom[797] = 12'h000;
rom[798] = 12'h00f;
rom[799] = 12'h00f;
rom[800] = 12'h00f;
rom[801] = 12'h00f;
rom[802] = 12'h00f;
rom[803] = 12'h00f;
rom[804] = 12'h000;
rom[805] = 12'h000;
rom[806] = 12'h000;
rom[807] = 12'h000;
rom[808] = 12'h000;
rom[809] = 12'h000;
rom[810] = 12'h007;
rom[811] = 12'h007;
rom[812] = 12'h000;
rom[813] = 12'h000;
rom[814] = 12'h000;
rom[815] = 12'h000;
rom[816] = 12'h000;
rom[817] = 12'h000;
rom[818] = 12'h000;
rom[819] = 12'h000;
rom[820] = 12'h000;
rom[821] = 12'h000;
rom[822] = 12'h000;
rom[823] = 12'h000;
rom[824] = 12'h00f;
rom[825] = 12'h00f;
rom[826] = 12'h00f;
rom[827] = 12'h00f;
rom[828] = 12'h00f;
rom[829] = 12'h00f;
rom[830] = 12'h000;
rom[831] = 12'h000;
rom[832] = 12'h000;
rom[833] = 12'h000;
rom[834] = 12'h007;
rom[835] = 12'h007;
rom[836] = 12'h000;
rom[837] = 12'h000;
rom[838] = 12'h007;
rom[839] = 12'h007;
rom[840] = 12'h000;
rom[841] = 12'h000;
rom[842] = 12'h000;
rom[843] = 12'h000;
rom[844] = 12'h000;
rom[845] = 12'h000;
rom[846] = 12'h000;
rom[847] = 12'h000;
rom[848] = 12'h000;
rom[849] = 12'h000;
rom[850] = 12'h00f;
rom[851] = 12'h00f;
rom[852] = 12'h00f;
rom[853] = 12'h00f;
rom[854] = 12'h00f;
rom[855] = 12'h00f;
rom[856] = 12'h000;
rom[857] = 12'h000;
rom[858] = 12'h000;
rom[859] = 12'h000;
rom[860] = 12'h007;
rom[861] = 12'h007;
rom[862] = 12'h000;
rom[863] = 12'h000;
rom[864] = 12'h007;
rom[865] = 12'h007;
rom[866] = 12'h000;
rom[867] = 12'h000;
rom[868] = 12'h000;
rom[869] = 12'h000;
rom[870] = 12'h000;
rom[871] = 12'h000;
rom[872] = 12'h000;
rom[873] = 12'h000;
rom[874] = 12'h000;
rom[875] = 12'h000;
rom[876] = 12'h00f;
rom[877] = 12'h00f;
rom[878] = 12'h00f;
rom[879] = 12'h00f;
rom[880] = 12'h00f;
rom[881] = 12'h00f;
rom[882] = 12'h000;
rom[883] = 12'h000;
rom[884] = 12'h000;
rom[885] = 12'h000;
rom[886] = 12'h000;
rom[887] = 12'h000;
rom[888] = 12'h007;
rom[889] = 12'h007;
rom[890] = 12'h000;
rom[891] = 12'h000;
rom[892] = 12'h000;
rom[893] = 12'h000;
rom[894] = 12'h000;
rom[895] = 12'h000;
rom[896] = 12'h000;
rom[897] = 12'h000;
rom[898] = 12'h000;
rom[899] = 12'h000;
rom[900] = 12'h000;
rom[901] = 12'h000;
rom[902] = 12'h00f;
rom[903] = 12'h00f;
rom[904] = 12'h00f;
rom[905] = 12'h00f;
rom[906] = 12'h00f;
rom[907] = 12'h00f;
rom[908] = 12'h000;
rom[909] = 12'h000;
rom[910] = 12'h000;
rom[911] = 12'h000;
rom[912] = 12'h000;
rom[913] = 12'h000;
rom[914] = 12'h007;
rom[915] = 12'h007;
rom[916] = 12'h000;
rom[917] = 12'h000;
rom[918] = 12'h000;
rom[919] = 12'h000;
rom[920] = 12'h000;
rom[921] = 12'h000;
rom[922] = 12'h000;
rom[923] = 12'h000;
rom[924] = 12'h000;
rom[925] = 12'h000;
rom[926] = 12'h000;
rom[927] = 12'h000;
rom[928] = 12'h00f;
rom[929] = 12'h00f;
rom[930] = 12'h00f;
rom[931] = 12'h00f;
rom[932] = 12'h00f;
rom[933] = 12'h00f;
rom[934] = 12'h000;
rom[935] = 12'h000;
rom[936] = 12'h000;
rom[937] = 12'h000;
rom[938] = 12'h007;
rom[939] = 12'h007;
rom[940] = 12'h000;
rom[941] = 12'h000;
rom[942] = 12'h007;
rom[943] = 12'h007;
rom[944] = 12'h000;
rom[945] = 12'h000;
rom[946] = 12'h000;
rom[947] = 12'h000;
rom[948] = 12'h000;
rom[949] = 12'h000;
rom[950] = 12'h000;
rom[951] = 12'h000;
rom[952] = 12'h000;
rom[953] = 12'h000;
rom[954] = 12'h00f;
rom[955] = 12'h00f;
rom[956] = 12'h00f;
rom[957] = 12'h00f;
rom[958] = 12'h00f;
rom[959] = 12'h00f;
rom[960] = 12'h000;
rom[961] = 12'h000;
rom[962] = 12'h000;
rom[963] = 12'h000;
rom[964] = 12'h007;
rom[965] = 12'h007;
rom[966] = 12'h000;
rom[967] = 12'h000;
rom[968] = 12'h007;
rom[969] = 12'h007;
rom[970] = 12'h000;
rom[971] = 12'h000;
rom[972] = 12'h000;
rom[973] = 12'h000;
rom[974] = 12'h000;
rom[975] = 12'h000;
rom[976] = 12'h000;
rom[977] = 12'h000;
rom[978] = 12'h000;
rom[979] = 12'h000;
rom[980] = 12'h00f;
rom[981] = 12'h00f;
rom[982] = 12'h00f;
rom[983] = 12'h00f;
rom[984] = 12'h00f;
rom[985] = 12'h00f;
rom[986] = 12'h000;
rom[987] = 12'h000;
rom[988] = 12'h000;
rom[989] = 12'h000;
rom[990] = 12'h000;
rom[991] = 12'h000;
rom[992] = 12'h007;
rom[993] = 12'h007;
rom[994] = 12'h000;
rom[995] = 12'h000;
rom[996] = 12'h00f;
rom[997] = 12'h00f;
rom[998] = 12'h00f;
rom[999] = 12'h00f;
rom[1000] = 12'h00f;
rom[1001] = 12'h00f;
rom[1002] = 12'h00f;
rom[1003] = 12'h00f;
rom[1004] = 12'h00f;
rom[1005] = 12'h00f;
rom[1006] = 12'h000;
rom[1007] = 12'h000;
rom[1008] = 12'h00f;
rom[1009] = 12'h00f;
rom[1010] = 12'h00f;
rom[1011] = 12'h00f;
rom[1012] = 12'h000;
rom[1013] = 12'h000;
rom[1014] = 12'h000;
rom[1015] = 12'h000;
rom[1016] = 12'h000;
rom[1017] = 12'h000;
rom[1018] = 12'h007;
rom[1019] = 12'h007;
rom[1020] = 12'h000;
rom[1021] = 12'h000;
rom[1022] = 12'h00f;
rom[1023] = 12'h00f;
rom[1024] = 12'h00f;
rom[1025] = 12'h00f;
rom[1026] = 12'h00f;
rom[1027] = 12'h00f;
rom[1028] = 12'h00f;
rom[1029] = 12'h00f;
rom[1030] = 12'h00f;
rom[1031] = 12'h00f;
rom[1032] = 12'h000;
rom[1033] = 12'h000;
rom[1034] = 12'h00f;
rom[1035] = 12'h00f;
rom[1036] = 12'h00f;
rom[1037] = 12'h00f;
rom[1038] = 12'h000;
rom[1039] = 12'h000;
rom[1040] = 12'h000;
rom[1041] = 12'h000;
rom[1042] = 12'h007;
rom[1043] = 12'h007;
rom[1044] = 12'h000;
rom[1045] = 12'h000;
rom[1046] = 12'h00f;
rom[1047] = 12'h00f;
rom[1048] = 12'h00f;
rom[1049] = 12'h00f;
rom[1050] = 12'h00f;
rom[1051] = 12'h00f;
rom[1052] = 12'h00f;
rom[1053] = 12'h00f;
rom[1054] = 12'h00f;
rom[1055] = 12'h00f;
rom[1056] = 12'h00f;
rom[1057] = 12'h00f;
rom[1058] = 12'h00f;
rom[1059] = 12'h00f;
rom[1060] = 12'h000;
rom[1061] = 12'h000;
rom[1062] = 12'h00f;
rom[1063] = 12'h00f;
rom[1064] = 12'h000;
rom[1065] = 12'h000;
rom[1066] = 12'h000;
rom[1067] = 12'h000;
rom[1068] = 12'h007;
rom[1069] = 12'h007;
rom[1070] = 12'h000;
rom[1071] = 12'h000;
rom[1072] = 12'h00f;
rom[1073] = 12'h00f;
rom[1074] = 12'h00f;
rom[1075] = 12'h00f;
rom[1076] = 12'h00f;
rom[1077] = 12'h00f;
rom[1078] = 12'h00f;
rom[1079] = 12'h00f;
rom[1080] = 12'h00f;
rom[1081] = 12'h00f;
rom[1082] = 12'h00f;
rom[1083] = 12'h00f;
rom[1084] = 12'h00f;
rom[1085] = 12'h00f;
rom[1086] = 12'h000;
rom[1087] = 12'h000;
rom[1088] = 12'h00f;
rom[1089] = 12'h00f;
rom[1090] = 12'h000;
rom[1091] = 12'h000;
rom[1092] = 12'h000;
rom[1093] = 12'h000;
rom[1094] = 12'h000;
rom[1095] = 12'h000;
rom[1096] = 12'h00f;
rom[1097] = 12'h00f;
rom[1098] = 12'h00f;
rom[1099] = 12'h00f;
rom[1100] = 12'h00f;
rom[1101] = 12'h00f;
rom[1102] = 12'h00f;
rom[1103] = 12'h00f;
rom[1104] = 12'h00f;
rom[1105] = 12'h00f;
rom[1106] = 12'h00f;
rom[1107] = 12'h00f;
rom[1108] = 12'h00f;
rom[1109] = 12'h00f;
rom[1110] = 12'h00f;
rom[1111] = 12'h00f;
rom[1112] = 12'h00f;
rom[1113] = 12'h00f;
rom[1114] = 12'h000;
rom[1115] = 12'h000;
rom[1116] = 12'h000;
rom[1117] = 12'h000;
rom[1118] = 12'h000;
rom[1119] = 12'h000;
rom[1120] = 12'h000;
rom[1121] = 12'h000;
rom[1122] = 12'h00f;
rom[1123] = 12'h00f;
rom[1124] = 12'h00f;
rom[1125] = 12'h00f;
rom[1126] = 12'h00f;
rom[1127] = 12'h00f;
rom[1128] = 12'h00f;
rom[1129] = 12'h00f;
rom[1130] = 12'h00f;
rom[1131] = 12'h00f;
rom[1132] = 12'h00f;
rom[1133] = 12'h00f;
rom[1134] = 12'h00f;
rom[1135] = 12'h00f;
rom[1136] = 12'h00f;
rom[1137] = 12'h00f;
rom[1138] = 12'h00f;
rom[1139] = 12'h00f;
rom[1140] = 12'h000;
rom[1141] = 12'h000;
rom[1142] = 12'h000;
rom[1143] = 12'h000;
rom[1144] = 12'h000;
rom[1145] = 12'h000;
rom[1146] = 12'h000;
rom[1147] = 12'h000;
rom[1148] = 12'h000;
rom[1149] = 12'h000;
rom[1150] = 12'h000;
rom[1151] = 12'h000;
rom[1152] = 12'h000;
rom[1153] = 12'h000;
rom[1154] = 12'h000;
rom[1155] = 12'h000;
rom[1156] = 12'h000;
rom[1157] = 12'h000;
rom[1158] = 12'h000;
rom[1159] = 12'h000;
rom[1160] = 12'h000;
rom[1161] = 12'h000;
rom[1162] = 12'h000;
rom[1163] = 12'h000;
rom[1164] = 12'h000;
rom[1165] = 12'h000;
rom[1166] = 12'h000;
rom[1167] = 12'h000;
rom[1168] = 12'h000;
rom[1169] = 12'h000;
rom[1170] = 12'h000;
rom[1171] = 12'h000;
rom[1172] = 12'h000;
rom[1173] = 12'h000;
rom[1174] = 12'h000;
rom[1175] = 12'h000;
rom[1176] = 12'h000;
rom[1177] = 12'h000;
rom[1178] = 12'h000;
rom[1179] = 12'h000;
rom[1180] = 12'h000;
rom[1181] = 12'h000;
rom[1182] = 12'h000;
rom[1183] = 12'h000;
rom[1184] = 12'h000;
rom[1185] = 12'h000;
rom[1186] = 12'h000;
rom[1187] = 12'h000;
rom[1188] = 12'h000;
rom[1189] = 12'h000;
rom[1190] = 12'h000;
rom[1191] = 12'h000;
rom[1192] = 12'h000;
rom[1193] = 12'h000;
rom[1194] = 12'h000;
rom[1195] = 12'h000;

  end
  endmodule

    module dash_rom (                       //четыре
  input  wire    [13:0]     addr,
  output wire    [11:0]     word
);

  logic [11:0] rom [(46 * 26)];

  assign word = rom[addr];

  initial begin
rom[0] = 12'h000;
rom[1] = 12'h000;
rom[2] = 12'h000;
rom[3] = 12'h000;
rom[4] = 12'h000;
rom[5] = 12'h000;
rom[6] = 12'h000;
rom[7] = 12'h000;
rom[8] = 12'h000;
rom[9] = 12'h000;
rom[10] = 12'h000;
rom[11] = 12'h000;
rom[12] = 12'h000;
rom[13] = 12'h000;
rom[14] = 12'h000;
rom[15] = 12'h000;
rom[16] = 12'h000;
rom[17] = 12'h000;
rom[18] = 12'h000;
rom[19] = 12'h000;
rom[20] = 12'h000;
rom[21] = 12'h000;
rom[22] = 12'h000;
rom[23] = 12'h000;
rom[24] = 12'h000;
rom[25] = 12'h000;
rom[26] = 12'h000;
rom[27] = 12'h000;
rom[28] = 12'h000;
rom[29] = 12'h000;
rom[30] = 12'h000;
rom[31] = 12'h000;
rom[32] = 12'h000;
rom[33] = 12'h000;
rom[34] = 12'h000;
rom[35] = 12'h000;
rom[36] = 12'h000;
rom[37] = 12'h000;
rom[38] = 12'h000;
rom[39] = 12'h000;
rom[40] = 12'h000;
rom[41] = 12'h000;
rom[42] = 12'h000;
rom[43] = 12'h000;
rom[44] = 12'h000;
rom[45] = 12'h000;
rom[46] = 12'h000;
rom[47] = 12'h000;
rom[48] = 12'h000;
rom[49] = 12'h000;
rom[50] = 12'h000;
rom[51] = 12'h000;
rom[52] = 12'h000;
rom[53] = 12'h000;
rom[54] = 12'h000;
rom[55] = 12'h000;
rom[56] = 12'h000;
rom[57] = 12'h000;
rom[58] = 12'h007;
rom[59] = 12'h007;
rom[60] = 12'h000;
rom[61] = 12'h000;
rom[62] = 12'h007;
rom[63] = 12'h007;
rom[64] = 12'h000;
rom[65] = 12'h000;
rom[66] = 12'h007;
rom[67] = 12'h007;
rom[68] = 12'h000;
rom[69] = 12'h000;
rom[70] = 12'h007;
rom[71] = 12'h007;
rom[72] = 12'h000;
rom[73] = 12'h000;
rom[74] = 12'h000;
rom[75] = 12'h000;
rom[76] = 12'h000;
rom[77] = 12'h000;
rom[78] = 12'h000;
rom[79] = 12'h000;
rom[80] = 12'h000;
rom[81] = 12'h000;
rom[82] = 12'h000;
rom[83] = 12'h000;
rom[84] = 12'h007;
rom[85] = 12'h007;
rom[86] = 12'h000;
rom[87] = 12'h000;
rom[88] = 12'h007;
rom[89] = 12'h007;
rom[90] = 12'h000;
rom[91] = 12'h000;
rom[92] = 12'h007;
rom[93] = 12'h007;
rom[94] = 12'h000;
rom[95] = 12'h000;
rom[96] = 12'h007;
rom[97] = 12'h007;
rom[98] = 12'h000;
rom[99] = 12'h000;
rom[100] = 12'h000;
rom[101] = 12'h000;
rom[102] = 12'h000;
rom[103] = 12'h000;
rom[104] = 12'h000;
rom[105] = 12'h000;
rom[106] = 12'h00f;
rom[107] = 12'h00f;
rom[108] = 12'h000;
rom[109] = 12'h000;
rom[110] = 12'h000;
rom[111] = 12'h000;
rom[112] = 12'h007;
rom[113] = 12'h007;
rom[114] = 12'h000;
rom[115] = 12'h000;
rom[116] = 12'h007;
rom[117] = 12'h007;
rom[118] = 12'h000;
rom[119] = 12'h000;
rom[120] = 12'h007;
rom[121] = 12'h007;
rom[122] = 12'h000;
rom[123] = 12'h000;
rom[124] = 12'h000;
rom[125] = 12'h000;
rom[126] = 12'h00f;
rom[127] = 12'h00f;
rom[128] = 12'h000;
rom[129] = 12'h000;
rom[130] = 12'h000;
rom[131] = 12'h000;
rom[132] = 12'h00f;
rom[133] = 12'h00f;
rom[134] = 12'h000;
rom[135] = 12'h000;
rom[136] = 12'h000;
rom[137] = 12'h000;
rom[138] = 12'h007;
rom[139] = 12'h007;
rom[140] = 12'h000;
rom[141] = 12'h000;
rom[142] = 12'h007;
rom[143] = 12'h007;
rom[144] = 12'h000;
rom[145] = 12'h000;
rom[146] = 12'h007;
rom[147] = 12'h007;
rom[148] = 12'h000;
rom[149] = 12'h000;
rom[150] = 12'h000;
rom[151] = 12'h000;
rom[152] = 12'h00f;
rom[153] = 12'h00f;
rom[154] = 12'h000;
rom[155] = 12'h000;
rom[156] = 12'h000;
rom[157] = 12'h000;
rom[158] = 12'h00f;
rom[159] = 12'h00f;
rom[160] = 12'h00f;
rom[161] = 12'h00f;
rom[162] = 12'h000;
rom[163] = 12'h000;
rom[164] = 12'h000;
rom[165] = 12'h000;
rom[166] = 12'h007;
rom[167] = 12'h007;
rom[168] = 12'h000;
rom[169] = 12'h000;
rom[170] = 12'h007;
rom[171] = 12'h007;
rom[172] = 12'h000;
rom[173] = 12'h000;
rom[174] = 12'h000;
rom[175] = 12'h000;
rom[176] = 12'h00f;
rom[177] = 12'h00f;
rom[178] = 12'h00f;
rom[179] = 12'h00f;
rom[180] = 12'h000;
rom[181] = 12'h000;
rom[182] = 12'h000;
rom[183] = 12'h000;
rom[184] = 12'h00f;
rom[185] = 12'h00f;
rom[186] = 12'h00f;
rom[187] = 12'h00f;
rom[188] = 12'h000;
rom[189] = 12'h000;
rom[190] = 12'h000;
rom[191] = 12'h000;
rom[192] = 12'h007;
rom[193] = 12'h007;
rom[194] = 12'h000;
rom[195] = 12'h000;
rom[196] = 12'h007;
rom[197] = 12'h007;
rom[198] = 12'h000;
rom[199] = 12'h000;
rom[200] = 12'h000;
rom[201] = 12'h000;
rom[202] = 12'h00f;
rom[203] = 12'h00f;
rom[204] = 12'h00f;
rom[205] = 12'h00f;
rom[206] = 12'h000;
rom[207] = 12'h000;
rom[208] = 12'h000;
rom[209] = 12'h000;
rom[210] = 12'h00f;
rom[211] = 12'h00f;
rom[212] = 12'h00f;
rom[213] = 12'h00f;
rom[214] = 12'h00f;
rom[215] = 12'h00f;
rom[216] = 12'h000;
rom[217] = 12'h000;
rom[218] = 12'h000;
rom[219] = 12'h000;
rom[220] = 12'h000;
rom[221] = 12'h000;
rom[222] = 12'h000;
rom[223] = 12'h000;
rom[224] = 12'h000;
rom[225] = 12'h000;
rom[226] = 12'h00f;
rom[227] = 12'h00f;
rom[228] = 12'h00f;
rom[229] = 12'h00f;
rom[230] = 12'h00f;
rom[231] = 12'h00f;
rom[232] = 12'h000;
rom[233] = 12'h000;
rom[234] = 12'h000;
rom[235] = 12'h000;
rom[236] = 12'h00f;
rom[237] = 12'h00f;
rom[238] = 12'h00f;
rom[239] = 12'h00f;
rom[240] = 12'h00f;
rom[241] = 12'h00f;
rom[242] = 12'h000;
rom[243] = 12'h000;
rom[244] = 12'h000;
rom[245] = 12'h000;
rom[246] = 12'h000;
rom[247] = 12'h000;
rom[248] = 12'h000;
rom[249] = 12'h000;
rom[250] = 12'h000;
rom[251] = 12'h000;
rom[252] = 12'h00f;
rom[253] = 12'h00f;
rom[254] = 12'h00f;
rom[255] = 12'h00f;
rom[256] = 12'h00f;
rom[257] = 12'h00f;
rom[258] = 12'h000;
rom[259] = 12'h000;
rom[260] = 12'h000;
rom[261] = 12'h000;
rom[262] = 12'h00f;
rom[263] = 12'h00f;
rom[264] = 12'h00f;
rom[265] = 12'h00f;
rom[266] = 12'h00f;
rom[267] = 12'h00f;
rom[268] = 12'h000;
rom[269] = 12'h000;
rom[270] = 12'h000;
rom[271] = 12'h000;
rom[272] = 12'h000;
rom[273] = 12'h000;
rom[274] = 12'h000;
rom[275] = 12'h000;
rom[276] = 12'h000;
rom[277] = 12'h000;
rom[278] = 12'h00f;
rom[279] = 12'h00f;
rom[280] = 12'h00f;
rom[281] = 12'h00f;
rom[282] = 12'h00f;
rom[283] = 12'h00f;
rom[284] = 12'h000;
rom[285] = 12'h000;
rom[286] = 12'h000;
rom[287] = 12'h000;
rom[288] = 12'h00f;
rom[289] = 12'h00f;
rom[290] = 12'h00f;
rom[291] = 12'h00f;
rom[292] = 12'h00f;
rom[293] = 12'h00f;
rom[294] = 12'h000;
rom[295] = 12'h000;
rom[296] = 12'h000;
rom[297] = 12'h000;
rom[298] = 12'h000;
rom[299] = 12'h000;
rom[300] = 12'h000;
rom[301] = 12'h000;
rom[302] = 12'h000;
rom[303] = 12'h000;
rom[304] = 12'h00f;
rom[305] = 12'h00f;
rom[306] = 12'h00f;
rom[307] = 12'h00f;
rom[308] = 12'h00f;
rom[309] = 12'h00f;
rom[310] = 12'h000;
rom[311] = 12'h000;
rom[312] = 12'h000;
rom[313] = 12'h000;
rom[314] = 12'h00f;
rom[315] = 12'h00f;
rom[316] = 12'h00f;
rom[317] = 12'h00f;
rom[318] = 12'h00f;
rom[319] = 12'h00f;
rom[320] = 12'h000;
rom[321] = 12'h000;
rom[322] = 12'h000;
rom[323] = 12'h000;
rom[324] = 12'h000;
rom[325] = 12'h000;
rom[326] = 12'h000;
rom[327] = 12'h000;
rom[328] = 12'h000;
rom[329] = 12'h000;
rom[330] = 12'h00f;
rom[331] = 12'h00f;
rom[332] = 12'h00f;
rom[333] = 12'h00f;
rom[334] = 12'h00f;
rom[335] = 12'h00f;
rom[336] = 12'h000;
rom[337] = 12'h000;
rom[338] = 12'h000;
rom[339] = 12'h000;
rom[340] = 12'h00f;
rom[341] = 12'h00f;
rom[342] = 12'h00f;
rom[343] = 12'h00f;
rom[344] = 12'h00f;
rom[345] = 12'h00f;
rom[346] = 12'h000;
rom[347] = 12'h000;
rom[348] = 12'h000;
rom[349] = 12'h000;
rom[350] = 12'h000;
rom[351] = 12'h000;
rom[352] = 12'h000;
rom[353] = 12'h000;
rom[354] = 12'h000;
rom[355] = 12'h000;
rom[356] = 12'h00f;
rom[357] = 12'h00f;
rom[358] = 12'h00f;
rom[359] = 12'h00f;
rom[360] = 12'h00f;
rom[361] = 12'h00f;
rom[362] = 12'h000;
rom[363] = 12'h000;
rom[364] = 12'h000;
rom[365] = 12'h000;
rom[366] = 12'h00f;
rom[367] = 12'h00f;
rom[368] = 12'h00f;
rom[369] = 12'h00f;
rom[370] = 12'h00f;
rom[371] = 12'h00f;
rom[372] = 12'h000;
rom[373] = 12'h000;
rom[374] = 12'h000;
rom[375] = 12'h000;
rom[376] = 12'h000;
rom[377] = 12'h000;
rom[378] = 12'h000;
rom[379] = 12'h000;
rom[380] = 12'h000;
rom[381] = 12'h000;
rom[382] = 12'h00f;
rom[383] = 12'h00f;
rom[384] = 12'h00f;
rom[385] = 12'h00f;
rom[386] = 12'h00f;
rom[387] = 12'h00f;
rom[388] = 12'h000;
rom[389] = 12'h000;
rom[390] = 12'h000;
rom[391] = 12'h000;
rom[392] = 12'h00f;
rom[393] = 12'h00f;
rom[394] = 12'h00f;
rom[395] = 12'h00f;
rom[396] = 12'h00f;
rom[397] = 12'h00f;
rom[398] = 12'h000;
rom[399] = 12'h000;
rom[400] = 12'h000;
rom[401] = 12'h000;
rom[402] = 12'h000;
rom[403] = 12'h000;
rom[404] = 12'h000;
rom[405] = 12'h000;
rom[406] = 12'h000;
rom[407] = 12'h000;
rom[408] = 12'h00f;
rom[409] = 12'h00f;
rom[410] = 12'h00f;
rom[411] = 12'h00f;
rom[412] = 12'h00f;
rom[413] = 12'h00f;
rom[414] = 12'h000;
rom[415] = 12'h000;
rom[416] = 12'h000;
rom[417] = 12'h000;
rom[418] = 12'h00f;
rom[419] = 12'h00f;
rom[420] = 12'h00f;
rom[421] = 12'h00f;
rom[422] = 12'h00f;
rom[423] = 12'h00f;
rom[424] = 12'h000;
rom[425] = 12'h000;
rom[426] = 12'h000;
rom[427] = 12'h000;
rom[428] = 12'h000;
rom[429] = 12'h000;
rom[430] = 12'h000;
rom[431] = 12'h000;
rom[432] = 12'h000;
rom[433] = 12'h000;
rom[434] = 12'h00f;
rom[435] = 12'h00f;
rom[436] = 12'h00f;
rom[437] = 12'h00f;
rom[438] = 12'h00f;
rom[439] = 12'h00f;
rom[440] = 12'h000;
rom[441] = 12'h000;
rom[442] = 12'h000;
rom[443] = 12'h000;
rom[444] = 12'h00f;
rom[445] = 12'h00f;
rom[446] = 12'h00f;
rom[447] = 12'h00f;
rom[448] = 12'h00f;
rom[449] = 12'h00f;
rom[450] = 12'h000;
rom[451] = 12'h000;
rom[452] = 12'h000;
rom[453] = 12'h000;
rom[454] = 12'h000;
rom[455] = 12'h000;
rom[456] = 12'h000;
rom[457] = 12'h000;
rom[458] = 12'h000;
rom[459] = 12'h000;
rom[460] = 12'h00f;
rom[461] = 12'h00f;
rom[462] = 12'h00f;
rom[463] = 12'h00f;
rom[464] = 12'h00f;
rom[465] = 12'h00f;
rom[466] = 12'h000;
rom[467] = 12'h000;
rom[468] = 12'h000;
rom[469] = 12'h000;
rom[470] = 12'h00f;
rom[471] = 12'h00f;
rom[472] = 12'h00f;
rom[473] = 12'h00f;
rom[474] = 12'h000;
rom[475] = 12'h000;
rom[476] = 12'h000;
rom[477] = 12'h000;
rom[478] = 12'h000;
rom[479] = 12'h000;
rom[480] = 12'h000;
rom[481] = 12'h000;
rom[482] = 12'h000;
rom[483] = 12'h000;
rom[484] = 12'h000;
rom[485] = 12'h000;
rom[486] = 12'h000;
rom[487] = 12'h000;
rom[488] = 12'h00f;
rom[489] = 12'h00f;
rom[490] = 12'h00f;
rom[491] = 12'h00f;
rom[492] = 12'h000;
rom[493] = 12'h000;
rom[494] = 12'h000;
rom[495] = 12'h000;
rom[496] = 12'h00f;
rom[497] = 12'h00f;
rom[498] = 12'h00f;
rom[499] = 12'h00f;
rom[500] = 12'h000;
rom[501] = 12'h000;
rom[502] = 12'h000;
rom[503] = 12'h000;
rom[504] = 12'h000;
rom[505] = 12'h000;
rom[506] = 12'h000;
rom[507] = 12'h000;
rom[508] = 12'h000;
rom[509] = 12'h000;
rom[510] = 12'h000;
rom[511] = 12'h000;
rom[512] = 12'h000;
rom[513] = 12'h000;
rom[514] = 12'h00f;
rom[515] = 12'h00f;
rom[516] = 12'h00f;
rom[517] = 12'h00f;
rom[518] = 12'h000;
rom[519] = 12'h000;
rom[520] = 12'h000;
rom[521] = 12'h000;
rom[522] = 12'h00f;
rom[523] = 12'h00f;
rom[524] = 12'h000;
rom[525] = 12'h000;
rom[526] = 12'h00f;
rom[527] = 12'h00f;
rom[528] = 12'h00f;
rom[529] = 12'h00f;
rom[530] = 12'h00f;
rom[531] = 12'h00f;
rom[532] = 12'h00f;
rom[533] = 12'h00f;
rom[534] = 12'h00f;
rom[535] = 12'h00f;
rom[536] = 12'h00f;
rom[537] = 12'h00f;
rom[538] = 12'h00f;
rom[539] = 12'h00f;
rom[540] = 12'h000;
rom[541] = 12'h000;
rom[542] = 12'h00f;
rom[543] = 12'h00f;
rom[544] = 12'h000;
rom[545] = 12'h000;
rom[546] = 12'h000;
rom[547] = 12'h000;
rom[548] = 12'h00f;
rom[549] = 12'h00f;
rom[550] = 12'h000;
rom[551] = 12'h000;
rom[552] = 12'h00f;
rom[553] = 12'h00f;
rom[554] = 12'h00f;
rom[555] = 12'h00f;
rom[556] = 12'h00f;
rom[557] = 12'h00f;
rom[558] = 12'h00f;
rom[559] = 12'h00f;
rom[560] = 12'h00f;
rom[561] = 12'h00f;
rom[562] = 12'h00f;
rom[563] = 12'h00f;
rom[564] = 12'h00f;
rom[565] = 12'h00f;
rom[566] = 12'h000;
rom[567] = 12'h000;
rom[568] = 12'h00f;
rom[569] = 12'h00f;
rom[570] = 12'h000;
rom[571] = 12'h000;
rom[572] = 12'h000;
rom[573] = 12'h000;
rom[574] = 12'h000;
rom[575] = 12'h000;
rom[576] = 12'h00f;
rom[577] = 12'h00f;
rom[578] = 12'h00f;
rom[579] = 12'h00f;
rom[580] = 12'h00f;
rom[581] = 12'h00f;
rom[582] = 12'h00f;
rom[583] = 12'h00f;
rom[584] = 12'h00f;
rom[585] = 12'h00f;
rom[586] = 12'h00f;
rom[587] = 12'h00f;
rom[588] = 12'h00f;
rom[589] = 12'h00f;
rom[590] = 12'h00f;
rom[591] = 12'h00f;
rom[592] = 12'h00f;
rom[593] = 12'h00f;
rom[594] = 12'h000;
rom[595] = 12'h000;
rom[596] = 12'h000;
rom[597] = 12'h000;
rom[598] = 12'h000;
rom[599] = 12'h000;
rom[600] = 12'h000;
rom[601] = 12'h000;
rom[602] = 12'h00f;
rom[603] = 12'h00f;
rom[604] = 12'h00f;
rom[605] = 12'h00f;
rom[606] = 12'h00f;
rom[607] = 12'h00f;
rom[608] = 12'h00f;
rom[609] = 12'h00f;
rom[610] = 12'h00f;
rom[611] = 12'h00f;
rom[612] = 12'h00f;
rom[613] = 12'h00f;
rom[614] = 12'h00f;
rom[615] = 12'h00f;
rom[616] = 12'h00f;
rom[617] = 12'h00f;
rom[618] = 12'h00f;
rom[619] = 12'h00f;
rom[620] = 12'h000;
rom[621] = 12'h000;
rom[622] = 12'h000;
rom[623] = 12'h000;
rom[624] = 12'h000;
rom[625] = 12'h000;
rom[626] = 12'h007;
rom[627] = 12'h007;
rom[628] = 12'h000;
rom[629] = 12'h000;
rom[630] = 12'h00f;
rom[631] = 12'h00f;
rom[632] = 12'h00f;
rom[633] = 12'h00f;
rom[634] = 12'h00f;
rom[635] = 12'h00f;
rom[636] = 12'h00f;
rom[637] = 12'h00f;
rom[638] = 12'h00f;
rom[639] = 12'h00f;
rom[640] = 12'h00f;
rom[641] = 12'h00f;
rom[642] = 12'h00f;
rom[643] = 12'h00f;
rom[644] = 12'h000;
rom[645] = 12'h000;
rom[646] = 12'h00f;
rom[647] = 12'h00f;
rom[648] = 12'h000;
rom[649] = 12'h000;
rom[650] = 12'h000;
rom[651] = 12'h000;
rom[652] = 12'h007;
rom[653] = 12'h007;
rom[654] = 12'h000;
rom[655] = 12'h000;
rom[656] = 12'h00f;
rom[657] = 12'h00f;
rom[658] = 12'h00f;
rom[659] = 12'h00f;
rom[660] = 12'h00f;
rom[661] = 12'h00f;
rom[662] = 12'h00f;
rom[663] = 12'h00f;
rom[664] = 12'h00f;
rom[665] = 12'h00f;
rom[666] = 12'h00f;
rom[667] = 12'h00f;
rom[668] = 12'h00f;
rom[669] = 12'h00f;
rom[670] = 12'h000;
rom[671] = 12'h000;
rom[672] = 12'h00f;
rom[673] = 12'h00f;
rom[674] = 12'h000;
rom[675] = 12'h000;
rom[676] = 12'h000;
rom[677] = 12'h000;
rom[678] = 12'h000;
rom[679] = 12'h000;
rom[680] = 12'h007;
rom[681] = 12'h007;
rom[682] = 12'h000;
rom[683] = 12'h000;
rom[684] = 12'h000;
rom[685] = 12'h000;
rom[686] = 12'h000;
rom[687] = 12'h000;
rom[688] = 12'h000;
rom[689] = 12'h000;
rom[690] = 12'h000;
rom[691] = 12'h000;
rom[692] = 12'h000;
rom[693] = 12'h000;
rom[694] = 12'h000;
rom[695] = 12'h000;
rom[696] = 12'h00f;
rom[697] = 12'h00f;
rom[698] = 12'h00f;
rom[699] = 12'h00f;
rom[700] = 12'h000;
rom[701] = 12'h000;
rom[702] = 12'h000;
rom[703] = 12'h000;
rom[704] = 12'h000;
rom[705] = 12'h000;
rom[706] = 12'h007;
rom[707] = 12'h007;
rom[708] = 12'h000;
rom[709] = 12'h000;
rom[710] = 12'h000;
rom[711] = 12'h000;
rom[712] = 12'h000;
rom[713] = 12'h000;
rom[714] = 12'h000;
rom[715] = 12'h000;
rom[716] = 12'h000;
rom[717] = 12'h000;
rom[718] = 12'h000;
rom[719] = 12'h000;
rom[720] = 12'h000;
rom[721] = 12'h000;
rom[722] = 12'h00f;
rom[723] = 12'h00f;
rom[724] = 12'h00f;
rom[725] = 12'h00f;
rom[726] = 12'h000;
rom[727] = 12'h000;
rom[728] = 12'h000;
rom[729] = 12'h000;
rom[730] = 12'h007;
rom[731] = 12'h007;
rom[732] = 12'h000;
rom[733] = 12'h000;
rom[734] = 12'h007;
rom[735] = 12'h007;
rom[736] = 12'h000;
rom[737] = 12'h000;
rom[738] = 12'h000;
rom[739] = 12'h000;
rom[740] = 12'h000;
rom[741] = 12'h000;
rom[742] = 12'h000;
rom[743] = 12'h000;
rom[744] = 12'h000;
rom[745] = 12'h000;
rom[746] = 12'h00f;
rom[747] = 12'h00f;
rom[748] = 12'h00f;
rom[749] = 12'h00f;
rom[750] = 12'h00f;
rom[751] = 12'h00f;
rom[752] = 12'h000;
rom[753] = 12'h000;
rom[754] = 12'h000;
rom[755] = 12'h000;
rom[756] = 12'h007;
rom[757] = 12'h007;
rom[758] = 12'h000;
rom[759] = 12'h000;
rom[760] = 12'h007;
rom[761] = 12'h007;
rom[762] = 12'h000;
rom[763] = 12'h000;
rom[764] = 12'h000;
rom[765] = 12'h000;
rom[766] = 12'h000;
rom[767] = 12'h000;
rom[768] = 12'h000;
rom[769] = 12'h000;
rom[770] = 12'h000;
rom[771] = 12'h000;
rom[772] = 12'h00f;
rom[773] = 12'h00f;
rom[774] = 12'h00f;
rom[775] = 12'h00f;
rom[776] = 12'h00f;
rom[777] = 12'h00f;
rom[778] = 12'h000;
rom[779] = 12'h000;
rom[780] = 12'h000;
rom[781] = 12'h000;
rom[782] = 12'h000;
rom[783] = 12'h000;
rom[784] = 12'h007;
rom[785] = 12'h007;
rom[786] = 12'h000;
rom[787] = 12'h000;
rom[788] = 12'h000;
rom[789] = 12'h000;
rom[790] = 12'h000;
rom[791] = 12'h000;
rom[792] = 12'h000;
rom[793] = 12'h000;
rom[794] = 12'h000;
rom[795] = 12'h000;
rom[796] = 12'h000;
rom[797] = 12'h000;
rom[798] = 12'h00f;
rom[799] = 12'h00f;
rom[800] = 12'h00f;
rom[801] = 12'h00f;
rom[802] = 12'h00f;
rom[803] = 12'h00f;
rom[804] = 12'h000;
rom[805] = 12'h000;
rom[806] = 12'h000;
rom[807] = 12'h000;
rom[808] = 12'h000;
rom[809] = 12'h000;
rom[810] = 12'h007;
rom[811] = 12'h007;
rom[812] = 12'h000;
rom[813] = 12'h000;
rom[814] = 12'h000;
rom[815] = 12'h000;
rom[816] = 12'h000;
rom[817] = 12'h000;
rom[818] = 12'h000;
rom[819] = 12'h000;
rom[820] = 12'h000;
rom[821] = 12'h000;
rom[822] = 12'h000;
rom[823] = 12'h000;
rom[824] = 12'h00f;
rom[825] = 12'h00f;
rom[826] = 12'h00f;
rom[827] = 12'h00f;
rom[828] = 12'h00f;
rom[829] = 12'h00f;
rom[830] = 12'h000;
rom[831] = 12'h000;
rom[832] = 12'h000;
rom[833] = 12'h000;
rom[834] = 12'h007;
rom[835] = 12'h007;
rom[836] = 12'h000;
rom[837] = 12'h000;
rom[838] = 12'h007;
rom[839] = 12'h007;
rom[840] = 12'h000;
rom[841] = 12'h000;
rom[842] = 12'h000;
rom[843] = 12'h000;
rom[844] = 12'h000;
rom[845] = 12'h000;
rom[846] = 12'h000;
rom[847] = 12'h000;
rom[848] = 12'h000;
rom[849] = 12'h000;
rom[850] = 12'h00f;
rom[851] = 12'h00f;
rom[852] = 12'h00f;
rom[853] = 12'h00f;
rom[854] = 12'h00f;
rom[855] = 12'h00f;
rom[856] = 12'h000;
rom[857] = 12'h000;
rom[858] = 12'h000;
rom[859] = 12'h000;
rom[860] = 12'h007;
rom[861] = 12'h007;
rom[862] = 12'h000;
rom[863] = 12'h000;
rom[864] = 12'h007;
rom[865] = 12'h007;
rom[866] = 12'h000;
rom[867] = 12'h000;
rom[868] = 12'h000;
rom[869] = 12'h000;
rom[870] = 12'h000;
rom[871] = 12'h000;
rom[872] = 12'h000;
rom[873] = 12'h000;
rom[874] = 12'h000;
rom[875] = 12'h000;
rom[876] = 12'h00f;
rom[877] = 12'h00f;
rom[878] = 12'h00f;
rom[879] = 12'h00f;
rom[880] = 12'h00f;
rom[881] = 12'h00f;
rom[882] = 12'h000;
rom[883] = 12'h000;
rom[884] = 12'h000;
rom[885] = 12'h000;
rom[886] = 12'h000;
rom[887] = 12'h000;
rom[888] = 12'h007;
rom[889] = 12'h007;
rom[890] = 12'h000;
rom[891] = 12'h000;
rom[892] = 12'h000;
rom[893] = 12'h000;
rom[894] = 12'h000;
rom[895] = 12'h000;
rom[896] = 12'h000;
rom[897] = 12'h000;
rom[898] = 12'h000;
rom[899] = 12'h000;
rom[900] = 12'h000;
rom[901] = 12'h000;
rom[902] = 12'h00f;
rom[903] = 12'h00f;
rom[904] = 12'h00f;
rom[905] = 12'h00f;
rom[906] = 12'h00f;
rom[907] = 12'h00f;
rom[908] = 12'h000;
rom[909] = 12'h000;
rom[910] = 12'h000;
rom[911] = 12'h000;
rom[912] = 12'h000;
rom[913] = 12'h000;
rom[914] = 12'h007;
rom[915] = 12'h007;
rom[916] = 12'h000;
rom[917] = 12'h000;
rom[918] = 12'h000;
rom[919] = 12'h000;
rom[920] = 12'h000;
rom[921] = 12'h000;
rom[922] = 12'h000;
rom[923] = 12'h000;
rom[924] = 12'h000;
rom[925] = 12'h000;
rom[926] = 12'h000;
rom[927] = 12'h000;
rom[928] = 12'h00f;
rom[929] = 12'h00f;
rom[930] = 12'h00f;
rom[931] = 12'h00f;
rom[932] = 12'h00f;
rom[933] = 12'h00f;
rom[934] = 12'h000;
rom[935] = 12'h000;
rom[936] = 12'h000;
rom[937] = 12'h000;
rom[938] = 12'h007;
rom[939] = 12'h007;
rom[940] = 12'h000;
rom[941] = 12'h000;
rom[942] = 12'h007;
rom[943] = 12'h007;
rom[944] = 12'h000;
rom[945] = 12'h000;
rom[946] = 12'h000;
rom[947] = 12'h000;
rom[948] = 12'h000;
rom[949] = 12'h000;
rom[950] = 12'h000;
rom[951] = 12'h000;
rom[952] = 12'h000;
rom[953] = 12'h000;
rom[954] = 12'h00f;
rom[955] = 12'h00f;
rom[956] = 12'h00f;
rom[957] = 12'h00f;
rom[958] = 12'h00f;
rom[959] = 12'h00f;
rom[960] = 12'h000;
rom[961] = 12'h000;
rom[962] = 12'h000;
rom[963] = 12'h000;
rom[964] = 12'h007;
rom[965] = 12'h007;
rom[966] = 12'h000;
rom[967] = 12'h000;
rom[968] = 12'h007;
rom[969] = 12'h007;
rom[970] = 12'h000;
rom[971] = 12'h000;
rom[972] = 12'h000;
rom[973] = 12'h000;
rom[974] = 12'h000;
rom[975] = 12'h000;
rom[976] = 12'h000;
rom[977] = 12'h000;
rom[978] = 12'h000;
rom[979] = 12'h000;
rom[980] = 12'h00f;
rom[981] = 12'h00f;
rom[982] = 12'h00f;
rom[983] = 12'h00f;
rom[984] = 12'h00f;
rom[985] = 12'h00f;
rom[986] = 12'h000;
rom[987] = 12'h000;
rom[988] = 12'h000;
rom[989] = 12'h000;
rom[990] = 12'h000;
rom[991] = 12'h000;
rom[992] = 12'h007;
rom[993] = 12'h007;
rom[994] = 12'h000;
rom[995] = 12'h000;
rom[996] = 12'h000;
rom[997] = 12'h000;
rom[998] = 12'h007;
rom[999] = 12'h007;
rom[1000] = 12'h000;
rom[1001] = 12'h000;
rom[1002] = 12'h007;
rom[1003] = 12'h007;
rom[1004] = 12'h000;
rom[1005] = 12'h000;
rom[1006] = 12'h000;
rom[1007] = 12'h000;
rom[1008] = 12'h00f;
rom[1009] = 12'h00f;
rom[1010] = 12'h00f;
rom[1011] = 12'h00f;
rom[1012] = 12'h000;
rom[1013] = 12'h000;
rom[1014] = 12'h000;
rom[1015] = 12'h000;
rom[1016] = 12'h000;
rom[1017] = 12'h000;
rom[1018] = 12'h007;
rom[1019] = 12'h007;
rom[1020] = 12'h000;
rom[1021] = 12'h000;
rom[1022] = 12'h000;
rom[1023] = 12'h000;
rom[1024] = 12'h007;
rom[1025] = 12'h007;
rom[1026] = 12'h000;
rom[1027] = 12'h000;
rom[1028] = 12'h007;
rom[1029] = 12'h007;
rom[1030] = 12'h000;
rom[1031] = 12'h000;
rom[1032] = 12'h000;
rom[1033] = 12'h000;
rom[1034] = 12'h00f;
rom[1035] = 12'h00f;
rom[1036] = 12'h00f;
rom[1037] = 12'h00f;
rom[1038] = 12'h000;
rom[1039] = 12'h000;
rom[1040] = 12'h000;
rom[1041] = 12'h000;
rom[1042] = 12'h007;
rom[1043] = 12'h007;
rom[1044] = 12'h000;
rom[1045] = 12'h000;
rom[1046] = 12'h000;
rom[1047] = 12'h000;
rom[1048] = 12'h007;
rom[1049] = 12'h007;
rom[1050] = 12'h000;
rom[1051] = 12'h000;
rom[1052] = 12'h007;
rom[1053] = 12'h007;
rom[1054] = 12'h000;
rom[1055] = 12'h000;
rom[1056] = 12'h007;
rom[1057] = 12'h007;
rom[1058] = 12'h000;
rom[1059] = 12'h000;
rom[1060] = 12'h000;
rom[1061] = 12'h000;
rom[1062] = 12'h00f;
rom[1063] = 12'h00f;
rom[1064] = 12'h000;
rom[1065] = 12'h000;
rom[1066] = 12'h000;
rom[1067] = 12'h000;
rom[1068] = 12'h007;
rom[1069] = 12'h007;
rom[1070] = 12'h000;
rom[1071] = 12'h000;
rom[1072] = 12'h000;
rom[1073] = 12'h000;
rom[1074] = 12'h007;
rom[1075] = 12'h007;
rom[1076] = 12'h000;
rom[1077] = 12'h000;
rom[1078] = 12'h007;
rom[1079] = 12'h007;
rom[1080] = 12'h000;
rom[1081] = 12'h000;
rom[1082] = 12'h007;
rom[1083] = 12'h007;
rom[1084] = 12'h000;
rom[1085] = 12'h000;
rom[1086] = 12'h000;
rom[1087] = 12'h000;
rom[1088] = 12'h00f;
rom[1089] = 12'h00f;
rom[1090] = 12'h000;
rom[1091] = 12'h000;
rom[1092] = 12'h000;
rom[1093] = 12'h000;
rom[1094] = 12'h000;
rom[1095] = 12'h000;
rom[1096] = 12'h000;
rom[1097] = 12'h000;
rom[1098] = 12'h007;
rom[1099] = 12'h007;
rom[1100] = 12'h000;
rom[1101] = 12'h000;
rom[1102] = 12'h007;
rom[1103] = 12'h007;
rom[1104] = 12'h000;
rom[1105] = 12'h000;
rom[1106] = 12'h007;
rom[1107] = 12'h007;
rom[1108] = 12'h000;
rom[1109] = 12'h000;
rom[1110] = 12'h007;
rom[1111] = 12'h007;
rom[1112] = 12'h000;
rom[1113] = 12'h000;
rom[1114] = 12'h000;
rom[1115] = 12'h000;
rom[1116] = 12'h000;
rom[1117] = 12'h000;
rom[1118] = 12'h000;
rom[1119] = 12'h000;
rom[1120] = 12'h000;
rom[1121] = 12'h000;
rom[1122] = 12'h000;
rom[1123] = 12'h000;
rom[1124] = 12'h007;
rom[1125] = 12'h007;
rom[1126] = 12'h000;
rom[1127] = 12'h000;
rom[1128] = 12'h007;
rom[1129] = 12'h007;
rom[1130] = 12'h000;
rom[1131] = 12'h000;
rom[1132] = 12'h007;
rom[1133] = 12'h007;
rom[1134] = 12'h000;
rom[1135] = 12'h000;
rom[1136] = 12'h007;
rom[1137] = 12'h007;
rom[1138] = 12'h000;
rom[1139] = 12'h000;
rom[1140] = 12'h000;
rom[1141] = 12'h000;
rom[1142] = 12'h000;
rom[1143] = 12'h000;
rom[1144] = 12'h000;
rom[1145] = 12'h000;
rom[1146] = 12'h000;
rom[1147] = 12'h000;
rom[1148] = 12'h000;
rom[1149] = 12'h000;
rom[1150] = 12'h000;
rom[1151] = 12'h000;
rom[1152] = 12'h000;
rom[1153] = 12'h000;
rom[1154] = 12'h000;
rom[1155] = 12'h000;
rom[1156] = 12'h000;
rom[1157] = 12'h000;
rom[1158] = 12'h000;
rom[1159] = 12'h000;
rom[1160] = 12'h000;
rom[1161] = 12'h000;
rom[1162] = 12'h000;
rom[1163] = 12'h000;
rom[1164] = 12'h000;
rom[1165] = 12'h000;
rom[1166] = 12'h000;
rom[1167] = 12'h000;
rom[1168] = 12'h000;
rom[1169] = 12'h000;
rom[1170] = 12'h000;
rom[1171] = 12'h000;
rom[1172] = 12'h000;
rom[1173] = 12'h000;
rom[1174] = 12'h000;
rom[1175] = 12'h000;
rom[1176] = 12'h000;
rom[1177] = 12'h000;
rom[1178] = 12'h000;
rom[1179] = 12'h000;
rom[1180] = 12'h000;
rom[1181] = 12'h000;
rom[1182] = 12'h000;
rom[1183] = 12'h000;
rom[1184] = 12'h000;
rom[1185] = 12'h000;
rom[1186] = 12'h000;
rom[1187] = 12'h000;
rom[1188] = 12'h000;
rom[1189] = 12'h000;
rom[1190] = 12'h000;
rom[1191] = 12'h000;
rom[1192] = 12'h000;
rom[1193] = 12'h000;
rom[1194] = 12'h000;
rom[1195] = 12'h000;
  end
  endmodule

    module dash_rom (                       //пять
  input  wire    [13:0]     addr,
  output wire    [11:0]     word
);

  logic [11:0] rom [(46 * 26)];

  assign word = rom[addr];

  initial begin
rom[0] = 12'h000;
rom[1] = 12'h000;
rom[2] = 12'h000;
rom[3] = 12'h000;
rom[4] = 12'h000;
rom[5] = 12'h000;
rom[6] = 12'h000;
rom[7] = 12'h000;
rom[8] = 12'h000;
rom[9] = 12'h000;
rom[10] = 12'h000;
rom[11] = 12'h000;
rom[12] = 12'h000;
rom[13] = 12'h000;
rom[14] = 12'h000;
rom[15] = 12'h000;
rom[16] = 12'h000;
rom[17] = 12'h000;
rom[18] = 12'h000;
rom[19] = 12'h000;
rom[20] = 12'h000;
rom[21] = 12'h000;
rom[22] = 12'h000;
rom[23] = 12'h000;
rom[24] = 12'h000;
rom[25] = 12'h000;
rom[26] = 12'h000;
rom[27] = 12'h000;
rom[28] = 12'h000;
rom[29] = 12'h000;
rom[30] = 12'h000;
rom[31] = 12'h000;
rom[32] = 12'h000;
rom[33] = 12'h000;
rom[34] = 12'h000;
rom[35] = 12'h000;
rom[36] = 12'h000;
rom[37] = 12'h000;
rom[38] = 12'h000;
rom[39] = 12'h000;
rom[40] = 12'h000;
rom[41] = 12'h000;
rom[42] = 12'h000;
rom[43] = 12'h000;
rom[44] = 12'h000;
rom[45] = 12'h000;
rom[46] = 12'h000;
rom[47] = 12'h000;
rom[48] = 12'h000;
rom[49] = 12'h000;
rom[50] = 12'h000;
rom[51] = 12'h000;
rom[52] = 12'h000;
rom[53] = 12'h000;
rom[54] = 12'h000;
rom[55] = 12'h000;
rom[56] = 12'h00f;
rom[57] = 12'h00f;
rom[58] = 12'h00f;
rom[59] = 12'h00f;
rom[60] = 12'h00f;
rom[61] = 12'h00f;
rom[62] = 12'h00f;
rom[63] = 12'h00f;
rom[64] = 12'h00f;
rom[65] = 12'h00f;
rom[66] = 12'h00f;
rom[67] = 12'h00f;
rom[68] = 12'h00f;
rom[69] = 12'h00f;
rom[70] = 12'h00f;
rom[71] = 12'h00f;
rom[72] = 12'h00f;
rom[73] = 12'h00f;
rom[74] = 12'h000;
rom[75] = 12'h000;
rom[76] = 12'h000;
rom[77] = 12'h000;
rom[78] = 12'h000;
rom[79] = 12'h000;
rom[80] = 12'h000;
rom[81] = 12'h000;
rom[82] = 12'h00f;
rom[83] = 12'h00f;
rom[84] = 12'h00f;
rom[85] = 12'h00f;
rom[86] = 12'h00f;
rom[87] = 12'h00f;
rom[88] = 12'h00f;
rom[89] = 12'h00f;
rom[90] = 12'h00f;
rom[91] = 12'h00f;
rom[92] = 12'h00f;
rom[93] = 12'h00f;
rom[94] = 12'h00f;
rom[95] = 12'h00f;
rom[96] = 12'h00f;
rom[97] = 12'h00f;
rom[98] = 12'h00f;
rom[99] = 12'h00f;
rom[100] = 12'h000;
rom[101] = 12'h000;
rom[102] = 12'h000;
rom[103] = 12'h000;
rom[104] = 12'h000;
rom[105] = 12'h000;
rom[106] = 12'h00f;
rom[107] = 12'h00f;
rom[108] = 12'h000;
rom[109] = 12'h000;
rom[110] = 12'h00f;
rom[111] = 12'h00f;
rom[112] = 12'h00f;
rom[113] = 12'h00f;
rom[114] = 12'h00f;
rom[115] = 12'h00f;
rom[116] = 12'h00f;
rom[117] = 12'h00f;
rom[118] = 12'h00f;
rom[119] = 12'h00f;
rom[120] = 12'h00f;
rom[121] = 12'h00f;
rom[122] = 12'h00f;
rom[123] = 12'h00f;
rom[124] = 12'h000;
rom[125] = 12'h000;
rom[126] = 12'h007;
rom[127] = 12'h007;
rom[128] = 12'h000;
rom[129] = 12'h000;
rom[130] = 12'h000;
rom[131] = 12'h000;
rom[132] = 12'h00f;
rom[133] = 12'h00f;
rom[134] = 12'h000;
rom[135] = 12'h000;
rom[136] = 12'h00f;
rom[137] = 12'h00f;
rom[138] = 12'h00f;
rom[139] = 12'h00f;
rom[140] = 12'h00f;
rom[141] = 12'h00f;
rom[142] = 12'h00f;
rom[143] = 12'h00f;
rom[144] = 12'h00f;
rom[145] = 12'h00f;
rom[146] = 12'h00f;
rom[147] = 12'h00f;
rom[148] = 12'h00f;
rom[149] = 12'h00f;
rom[150] = 12'h000;
rom[151] = 12'h000;
rom[152] = 12'h007;
rom[153] = 12'h007;
rom[154] = 12'h000;
rom[155] = 12'h000;
rom[156] = 12'h000;
rom[157] = 12'h000;
rom[158] = 12'h00f;
rom[159] = 12'h00f;
rom[160] = 12'h00f;
rom[161] = 12'h00f;
rom[162] = 12'h000;
rom[163] = 12'h000;
rom[164] = 12'h00f;
rom[165] = 12'h00f;
rom[166] = 12'h00f;
rom[167] = 12'h00f;
rom[168] = 12'h00f;
rom[169] = 12'h00f;
rom[170] = 12'h00f;
rom[171] = 12'h00f;
rom[172] = 12'h00f;
rom[173] = 12'h00f;
rom[174] = 12'h000;
rom[175] = 12'h000;
rom[176] = 12'h007;
rom[177] = 12'h007;
rom[178] = 12'h000;
rom[179] = 12'h000;
rom[180] = 12'h000;
rom[181] = 12'h000;
rom[182] = 12'h000;
rom[183] = 12'h000;
rom[184] = 12'h00f;
rom[185] = 12'h00f;
rom[186] = 12'h00f;
rom[187] = 12'h00f;
rom[188] = 12'h000;
rom[189] = 12'h000;
rom[190] = 12'h00f;
rom[191] = 12'h00f;
rom[192] = 12'h00f;
rom[193] = 12'h00f;
rom[194] = 12'h00f;
rom[195] = 12'h00f;
rom[196] = 12'h00f;
rom[197] = 12'h00f;
rom[198] = 12'h00f;
rom[199] = 12'h00f;
rom[200] = 12'h000;
rom[201] = 12'h000;
rom[202] = 12'h007;
rom[203] = 12'h007;
rom[204] = 12'h000;
rom[205] = 12'h000;
rom[206] = 12'h000;
rom[207] = 12'h000;
rom[208] = 12'h000;
rom[209] = 12'h000;
rom[210] = 12'h00f;
rom[211] = 12'h00f;
rom[212] = 12'h00f;
rom[213] = 12'h00f;
rom[214] = 12'h00f;
rom[215] = 12'h00f;
rom[216] = 12'h000;
rom[217] = 12'h000;
rom[218] = 12'h000;
rom[219] = 12'h000;
rom[220] = 12'h000;
rom[221] = 12'h000;
rom[222] = 12'h000;
rom[223] = 12'h000;
rom[224] = 12'h000;
rom[225] = 12'h000;
rom[226] = 12'h007;
rom[227] = 12'h007;
rom[228] = 12'h000;
rom[229] = 12'h000;
rom[230] = 12'h007;
rom[231] = 12'h007;
rom[232] = 12'h000;
rom[233] = 12'h000;
rom[234] = 12'h000;
rom[235] = 12'h000;
rom[236] = 12'h00f;
rom[237] = 12'h00f;
rom[238] = 12'h00f;
rom[239] = 12'h00f;
rom[240] = 12'h00f;
rom[241] = 12'h00f;
rom[242] = 12'h000;
rom[243] = 12'h000;
rom[244] = 12'h000;
rom[245] = 12'h000;
rom[246] = 12'h000;
rom[247] = 12'h000;
rom[248] = 12'h000;
rom[249] = 12'h000;
rom[250] = 12'h000;
rom[251] = 12'h000;
rom[252] = 12'h007;
rom[253] = 12'h007;
rom[254] = 12'h000;
rom[255] = 12'h000;
rom[256] = 12'h007;
rom[257] = 12'h007;
rom[258] = 12'h000;
rom[259] = 12'h000;
rom[260] = 12'h000;
rom[261] = 12'h000;
rom[262] = 12'h00f;
rom[263] = 12'h00f;
rom[264] = 12'h00f;
rom[265] = 12'h00f;
rom[266] = 12'h00f;
rom[267] = 12'h00f;
rom[268] = 12'h000;
rom[269] = 12'h000;
rom[270] = 12'h000;
rom[271] = 12'h000;
rom[272] = 12'h000;
rom[273] = 12'h000;
rom[274] = 12'h000;
rom[275] = 12'h000;
rom[276] = 12'h000;
rom[277] = 12'h000;
rom[278] = 12'h000;
rom[279] = 12'h000;
rom[280] = 12'h007;
rom[281] = 12'h007;
rom[282] = 12'h000;
rom[283] = 12'h000;
rom[284] = 12'h000;
rom[285] = 12'h000;
rom[286] = 12'h000;
rom[287] = 12'h000;
rom[288] = 12'h00f;
rom[289] = 12'h00f;
rom[290] = 12'h00f;
rom[291] = 12'h00f;
rom[292] = 12'h00f;
rom[293] = 12'h00f;
rom[294] = 12'h000;
rom[295] = 12'h000;
rom[296] = 12'h000;
rom[297] = 12'h000;
rom[298] = 12'h000;
rom[299] = 12'h000;
rom[300] = 12'h000;
rom[301] = 12'h000;
rom[302] = 12'h000;
rom[303] = 12'h000;
rom[304] = 12'h000;
rom[305] = 12'h000;
rom[306] = 12'h007;
rom[307] = 12'h007;
rom[308] = 12'h000;
rom[309] = 12'h000;
rom[310] = 12'h000;
rom[311] = 12'h000;
rom[312] = 12'h000;
rom[313] = 12'h000;
rom[314] = 12'h00f;
rom[315] = 12'h00f;
rom[316] = 12'h00f;
rom[317] = 12'h00f;
rom[318] = 12'h00f;
rom[319] = 12'h00f;
rom[320] = 12'h000;
rom[321] = 12'h000;
rom[322] = 12'h000;
rom[323] = 12'h000;
rom[324] = 12'h000;
rom[325] = 12'h000;
rom[326] = 12'h000;
rom[327] = 12'h000;
rom[328] = 12'h000;
rom[329] = 12'h000;
rom[330] = 12'h007;
rom[331] = 12'h007;
rom[332] = 12'h000;
rom[333] = 12'h000;
rom[334] = 12'h007;
rom[335] = 12'h007;
rom[336] = 12'h000;
rom[337] = 12'h000;
rom[338] = 12'h000;
rom[339] = 12'h000;
rom[340] = 12'h00f;
rom[341] = 12'h00f;
rom[342] = 12'h00f;
rom[343] = 12'h00f;
rom[344] = 12'h00f;
rom[345] = 12'h00f;
rom[346] = 12'h000;
rom[347] = 12'h000;
rom[348] = 12'h000;
rom[349] = 12'h000;
rom[350] = 12'h000;
rom[351] = 12'h000;
rom[352] = 12'h000;
rom[353] = 12'h000;
rom[354] = 12'h000;
rom[355] = 12'h000;
rom[356] = 12'h007;
rom[357] = 12'h007;
rom[358] = 12'h000;
rom[359] = 12'h000;
rom[360] = 12'h007;
rom[361] = 12'h007;
rom[362] = 12'h000;
rom[363] = 12'h000;
rom[364] = 12'h000;
rom[365] = 12'h000;
rom[366] = 12'h00f;
rom[367] = 12'h00f;
rom[368] = 12'h00f;
rom[369] = 12'h00f;
rom[370] = 12'h00f;
rom[371] = 12'h00f;
rom[372] = 12'h000;
rom[373] = 12'h000;
rom[374] = 12'h000;
rom[375] = 12'h000;
rom[376] = 12'h000;
rom[377] = 12'h000;
rom[378] = 12'h000;
rom[379] = 12'h000;
rom[380] = 12'h000;
rom[381] = 12'h000;
rom[382] = 12'h000;
rom[383] = 12'h000;
rom[384] = 12'h007;
rom[385] = 12'h007;
rom[386] = 12'h000;
rom[387] = 12'h000;
rom[388] = 12'h000;
rom[389] = 12'h000;
rom[390] = 12'h000;
rom[391] = 12'h000;
rom[392] = 12'h00f;
rom[393] = 12'h00f;
rom[394] = 12'h00f;
rom[395] = 12'h00f;
rom[396] = 12'h00f;
rom[397] = 12'h00f;
rom[398] = 12'h000;
rom[399] = 12'h000;
rom[400] = 12'h000;
rom[401] = 12'h000;
rom[402] = 12'h000;
rom[403] = 12'h000;
rom[404] = 12'h000;
rom[405] = 12'h000;
rom[406] = 12'h000;
rom[407] = 12'h000;
rom[408] = 12'h000;
rom[409] = 12'h000;
rom[410] = 12'h007;
rom[411] = 12'h007;
rom[412] = 12'h000;
rom[413] = 12'h000;
rom[414] = 12'h000;
rom[415] = 12'h000;
rom[416] = 12'h000;
rom[417] = 12'h000;
rom[418] = 12'h00f;
rom[419] = 12'h00f;
rom[420] = 12'h00f;
rom[421] = 12'h00f;
rom[422] = 12'h00f;
rom[423] = 12'h00f;
rom[424] = 12'h000;
rom[425] = 12'h000;
rom[426] = 12'h000;
rom[427] = 12'h000;
rom[428] = 12'h000;
rom[429] = 12'h000;
rom[430] = 12'h000;
rom[431] = 12'h000;
rom[432] = 12'h000;
rom[433] = 12'h000;
rom[434] = 12'h007;
rom[435] = 12'h007;
rom[436] = 12'h000;
rom[437] = 12'h000;
rom[438] = 12'h007;
rom[439] = 12'h007;
rom[440] = 12'h000;
rom[441] = 12'h000;
rom[442] = 12'h000;
rom[443] = 12'h000;
rom[444] = 12'h00f;
rom[445] = 12'h00f;
rom[446] = 12'h00f;
rom[447] = 12'h00f;
rom[448] = 12'h00f;
rom[449] = 12'h00f;
rom[450] = 12'h000;
rom[451] = 12'h000;
rom[452] = 12'h000;
rom[453] = 12'h000;
rom[454] = 12'h000;
rom[455] = 12'h000;
rom[456] = 12'h000;
rom[457] = 12'h000;
rom[458] = 12'h000;
rom[459] = 12'h000;
rom[460] = 12'h007;
rom[461] = 12'h007;
rom[462] = 12'h000;
rom[463] = 12'h000;
rom[464] = 12'h007;
rom[465] = 12'h007;
rom[466] = 12'h000;
rom[467] = 12'h000;
rom[468] = 12'h000;
rom[469] = 12'h000;
rom[470] = 12'h00f;
rom[471] = 12'h00f;
rom[472] = 12'h00f;
rom[473] = 12'h00f;
rom[474] = 12'h000;
rom[475] = 12'h000;
rom[476] = 12'h000;
rom[477] = 12'h000;
rom[478] = 12'h000;
rom[479] = 12'h000;
rom[480] = 12'h000;
rom[481] = 12'h000;
rom[482] = 12'h000;
rom[483] = 12'h000;
rom[484] = 12'h000;
rom[485] = 12'h000;
rom[486] = 12'h000;
rom[487] = 12'h000;
rom[488] = 12'h007;
rom[489] = 12'h007;
rom[490] = 12'h000;
rom[491] = 12'h000;
rom[492] = 12'h000;
rom[493] = 12'h000;
rom[494] = 12'h000;
rom[495] = 12'h000;
rom[496] = 12'h00f;
rom[497] = 12'h00f;
rom[498] = 12'h00f;
rom[499] = 12'h00f;
rom[500] = 12'h000;
rom[501] = 12'h000;
rom[502] = 12'h000;
rom[503] = 12'h000;
rom[504] = 12'h000;
rom[505] = 12'h000;
rom[506] = 12'h000;
rom[507] = 12'h000;
rom[508] = 12'h000;
rom[509] = 12'h000;
rom[510] = 12'h000;
rom[511] = 12'h000;
rom[512] = 12'h000;
rom[513] = 12'h000;
rom[514] = 12'h007;
rom[515] = 12'h007;
rom[516] = 12'h000;
rom[517] = 12'h000;
rom[518] = 12'h000;
rom[519] = 12'h000;
rom[520] = 12'h000;
rom[521] = 12'h000;
rom[522] = 12'h00f;
rom[523] = 12'h00f;
rom[524] = 12'h000;
rom[525] = 12'h000;
rom[526] = 12'h00f;
rom[527] = 12'h00f;
rom[528] = 12'h00f;
rom[529] = 12'h00f;
rom[530] = 12'h00f;
rom[531] = 12'h00f;
rom[532] = 12'h00f;
rom[533] = 12'h00f;
rom[534] = 12'h00f;
rom[535] = 12'h00f;
rom[536] = 12'h00f;
rom[537] = 12'h00f;
rom[538] = 12'h00f;
rom[539] = 12'h00f;
rom[540] = 12'h000;
rom[541] = 12'h000;
rom[542] = 12'h007;
rom[543] = 12'h007;
rom[544] = 12'h000;
rom[545] = 12'h000;
rom[546] = 12'h000;
rom[547] = 12'h000;
rom[548] = 12'h00f;
rom[549] = 12'h00f;
rom[550] = 12'h000;
rom[551] = 12'h000;
rom[552] = 12'h00f;
rom[553] = 12'h00f;
rom[554] = 12'h00f;
rom[555] = 12'h00f;
rom[556] = 12'h00f;
rom[557] = 12'h00f;
rom[558] = 12'h00f;
rom[559] = 12'h00f;
rom[560] = 12'h00f;
rom[561] = 12'h00f;
rom[562] = 12'h00f;
rom[563] = 12'h00f;
rom[564] = 12'h00f;
rom[565] = 12'h00f;
rom[566] = 12'h000;
rom[567] = 12'h000;
rom[568] = 12'h007;
rom[569] = 12'h007;
rom[570] = 12'h000;
rom[571] = 12'h000;
rom[572] = 12'h000;
rom[573] = 12'h000;
rom[574] = 12'h000;
rom[575] = 12'h000;
rom[576] = 12'h00f;
rom[577] = 12'h00f;
rom[578] = 12'h00f;
rom[579] = 12'h00f;
rom[580] = 12'h00f;
rom[581] = 12'h00f;
rom[582] = 12'h00f;
rom[583] = 12'h00f;
rom[584] = 12'h00f;
rom[585] = 12'h00f;
rom[586] = 12'h00f;
rom[587] = 12'h00f;
rom[588] = 12'h00f;
rom[589] = 12'h00f;
rom[590] = 12'h00f;
rom[591] = 12'h00f;
rom[592] = 12'h00f;
rom[593] = 12'h00f;
rom[594] = 12'h000;
rom[595] = 12'h000;
rom[596] = 12'h000;
rom[597] = 12'h000;
rom[598] = 12'h000;
rom[599] = 12'h000;
rom[600] = 12'h000;
rom[601] = 12'h000;
rom[602] = 12'h00f;
rom[603] = 12'h00f;
rom[604] = 12'h00f;
rom[605] = 12'h00f;
rom[606] = 12'h00f;
rom[607] = 12'h00f;
rom[608] = 12'h00f;
rom[609] = 12'h00f;
rom[610] = 12'h00f;
rom[611] = 12'h00f;
rom[612] = 12'h00f;
rom[613] = 12'h00f;
rom[614] = 12'h00f;
rom[615] = 12'h00f;
rom[616] = 12'h00f;
rom[617] = 12'h00f;
rom[618] = 12'h00f;
rom[619] = 12'h00f;
rom[620] = 12'h000;
rom[621] = 12'h000;
rom[622] = 12'h000;
rom[623] = 12'h000;
rom[624] = 12'h000;
rom[625] = 12'h000;
rom[626] = 12'h007;
rom[627] = 12'h007;
rom[628] = 12'h000;
rom[629] = 12'h000;
rom[630] = 12'h00f;
rom[631] = 12'h00f;
rom[632] = 12'h00f;
rom[633] = 12'h00f;
rom[634] = 12'h00f;
rom[635] = 12'h00f;
rom[636] = 12'h00f;
rom[637] = 12'h00f;
rom[638] = 12'h00f;
rom[639] = 12'h00f;
rom[640] = 12'h00f;
rom[641] = 12'h00f;
rom[642] = 12'h00f;
rom[643] = 12'h00f;
rom[644] = 12'h000;
rom[645] = 12'h000;
rom[646] = 12'h00f;
rom[647] = 12'h00f;
rom[648] = 12'h000;
rom[649] = 12'h000;
rom[650] = 12'h000;
rom[651] = 12'h000;
rom[652] = 12'h007;
rom[653] = 12'h007;
rom[654] = 12'h000;
rom[655] = 12'h000;
rom[656] = 12'h00f;
rom[657] = 12'h00f;
rom[658] = 12'h00f;
rom[659] = 12'h00f;
rom[660] = 12'h00f;
rom[661] = 12'h00f;
rom[662] = 12'h00f;
rom[663] = 12'h00f;
rom[664] = 12'h00f;
rom[665] = 12'h00f;
rom[666] = 12'h00f;
rom[667] = 12'h00f;
rom[668] = 12'h00f;
rom[669] = 12'h00f;
rom[670] = 12'h000;
rom[671] = 12'h000;
rom[672] = 12'h00f;
rom[673] = 12'h00f;
rom[674] = 12'h000;
rom[675] = 12'h000;
rom[676] = 12'h000;
rom[677] = 12'h000;
rom[678] = 12'h000;
rom[679] = 12'h000;
rom[680] = 12'h007;
rom[681] = 12'h007;
rom[682] = 12'h000;
rom[683] = 12'h000;
rom[684] = 12'h000;
rom[685] = 12'h000;
rom[686] = 12'h000;
rom[687] = 12'h000;
rom[688] = 12'h000;
rom[689] = 12'h000;
rom[690] = 12'h000;
rom[691] = 12'h000;
rom[692] = 12'h000;
rom[693] = 12'h000;
rom[694] = 12'h000;
rom[695] = 12'h000;
rom[696] = 12'h00f;
rom[697] = 12'h00f;
rom[698] = 12'h00f;
rom[699] = 12'h00f;
rom[700] = 12'h000;
rom[701] = 12'h000;
rom[702] = 12'h000;
rom[703] = 12'h000;
rom[704] = 12'h000;
rom[705] = 12'h000;
rom[706] = 12'h007;
rom[707] = 12'h007;
rom[708] = 12'h000;
rom[709] = 12'h000;
rom[710] = 12'h000;
rom[711] = 12'h000;
rom[712] = 12'h000;
rom[713] = 12'h000;
rom[714] = 12'h000;
rom[715] = 12'h000;
rom[716] = 12'h000;
rom[717] = 12'h000;
rom[718] = 12'h000;
rom[719] = 12'h000;
rom[720] = 12'h000;
rom[721] = 12'h000;
rom[722] = 12'h00f;
rom[723] = 12'h00f;
rom[724] = 12'h00f;
rom[725] = 12'h00f;
rom[726] = 12'h000;
rom[727] = 12'h000;
rom[728] = 12'h000;
rom[729] = 12'h000;
rom[730] = 12'h007;
rom[731] = 12'h007;
rom[732] = 12'h000;
rom[733] = 12'h000;
rom[734] = 12'h007;
rom[735] = 12'h007;
rom[736] = 12'h000;
rom[737] = 12'h000;
rom[738] = 12'h000;
rom[739] = 12'h000;
rom[740] = 12'h000;
rom[741] = 12'h000;
rom[742] = 12'h000;
rom[743] = 12'h000;
rom[744] = 12'h000;
rom[745] = 12'h000;
rom[746] = 12'h00f;
rom[747] = 12'h00f;
rom[748] = 12'h00f;
rom[749] = 12'h00f;
rom[750] = 12'h00f;
rom[751] = 12'h00f;
rom[752] = 12'h000;
rom[753] = 12'h000;
rom[754] = 12'h000;
rom[755] = 12'h000;
rom[756] = 12'h007;
rom[757] = 12'h007;
rom[758] = 12'h000;
rom[759] = 12'h000;
rom[760] = 12'h007;
rom[761] = 12'h007;
rom[762] = 12'h000;
rom[763] = 12'h000;
rom[764] = 12'h000;
rom[765] = 12'h000;
rom[766] = 12'h000;
rom[767] = 12'h000;
rom[768] = 12'h000;
rom[769] = 12'h000;
rom[770] = 12'h000;
rom[771] = 12'h000;
rom[772] = 12'h00f;
rom[773] = 12'h00f;
rom[774] = 12'h00f;
rom[775] = 12'h00f;
rom[776] = 12'h00f;
rom[777] = 12'h00f;
rom[778] = 12'h000;
rom[779] = 12'h000;
rom[780] = 12'h000;
rom[781] = 12'h000;
rom[782] = 12'h000;
rom[783] = 12'h000;
rom[784] = 12'h007;
rom[785] = 12'h007;
rom[786] = 12'h000;
rom[787] = 12'h000;
rom[788] = 12'h000;
rom[789] = 12'h000;
rom[790] = 12'h000;
rom[791] = 12'h000;
rom[792] = 12'h000;
rom[793] = 12'h000;
rom[794] = 12'h000;
rom[795] = 12'h000;
rom[796] = 12'h000;
rom[797] = 12'h000;
rom[798] = 12'h00f;
rom[799] = 12'h00f;
rom[800] = 12'h00f;
rom[801] = 12'h00f;
rom[802] = 12'h00f;
rom[803] = 12'h00f;
rom[804] = 12'h000;
rom[805] = 12'h000;
rom[806] = 12'h000;
rom[807] = 12'h000;
rom[808] = 12'h000;
rom[809] = 12'h000;
rom[810] = 12'h007;
rom[811] = 12'h007;
rom[812] = 12'h000;
rom[813] = 12'h000;
rom[814] = 12'h000;
rom[815] = 12'h000;
rom[816] = 12'h000;
rom[817] = 12'h000;
rom[818] = 12'h000;
rom[819] = 12'h000;
rom[820] = 12'h000;
rom[821] = 12'h000;
rom[822] = 12'h000;
rom[823] = 12'h000;
rom[824] = 12'h00f;
rom[825] = 12'h00f;
rom[826] = 12'h00f;
rom[827] = 12'h00f;
rom[828] = 12'h00f;
rom[829] = 12'h00f;
rom[830] = 12'h000;
rom[831] = 12'h000;
rom[832] = 12'h000;
rom[833] = 12'h000;
rom[834] = 12'h007;
rom[835] = 12'h007;
rom[836] = 12'h000;
rom[837] = 12'h000;
rom[838] = 12'h007;
rom[839] = 12'h007;
rom[840] = 12'h000;
rom[841] = 12'h000;
rom[842] = 12'h000;
rom[843] = 12'h000;
rom[844] = 12'h000;
rom[845] = 12'h000;
rom[846] = 12'h000;
rom[847] = 12'h000;
rom[848] = 12'h000;
rom[849] = 12'h000;
rom[850] = 12'h00f;
rom[851] = 12'h00f;
rom[852] = 12'h00f;
rom[853] = 12'h00f;
rom[854] = 12'h00f;
rom[855] = 12'h00f;
rom[856] = 12'h000;
rom[857] = 12'h000;
rom[858] = 12'h000;
rom[859] = 12'h000;
rom[860] = 12'h007;
rom[861] = 12'h007;
rom[862] = 12'h000;
rom[863] = 12'h000;
rom[864] = 12'h007;
rom[865] = 12'h007;
rom[866] = 12'h000;
rom[867] = 12'h000;
rom[868] = 12'h000;
rom[869] = 12'h000;
rom[870] = 12'h000;
rom[871] = 12'h000;
rom[872] = 12'h000;
rom[873] = 12'h000;
rom[874] = 12'h000;
rom[875] = 12'h000;
rom[876] = 12'h00f;
rom[877] = 12'h00f;
rom[878] = 12'h00f;
rom[879] = 12'h00f;
rom[880] = 12'h00f;
rom[881] = 12'h00f;
rom[882] = 12'h000;
rom[883] = 12'h000;
rom[884] = 12'h000;
rom[885] = 12'h000;
rom[886] = 12'h000;
rom[887] = 12'h000;
rom[888] = 12'h007;
rom[889] = 12'h007;
rom[890] = 12'h000;
rom[891] = 12'h000;
rom[892] = 12'h000;
rom[893] = 12'h000;
rom[894] = 12'h000;
rom[895] = 12'h000;
rom[896] = 12'h000;
rom[897] = 12'h000;
rom[898] = 12'h000;
rom[899] = 12'h000;
rom[900] = 12'h000;
rom[901] = 12'h000;
rom[902] = 12'h00f;
rom[903] = 12'h00f;
rom[904] = 12'h00f;
rom[905] = 12'h00f;
rom[906] = 12'h00f;
rom[907] = 12'h00f;
rom[908] = 12'h000;
rom[909] = 12'h000;
rom[910] = 12'h000;
rom[911] = 12'h000;
rom[912] = 12'h000;
rom[913] = 12'h000;
rom[914] = 12'h007;
rom[915] = 12'h007;
rom[916] = 12'h000;
rom[917] = 12'h000;
rom[918] = 12'h000;
rom[919] = 12'h000;
rom[920] = 12'h000;
rom[921] = 12'h000;
rom[922] = 12'h000;
rom[923] = 12'h000;
rom[924] = 12'h000;
rom[925] = 12'h000;
rom[926] = 12'h000;
rom[927] = 12'h000;
rom[928] = 12'h00f;
rom[929] = 12'h00f;
rom[930] = 12'h00f;
rom[931] = 12'h00f;
rom[932] = 12'h00f;
rom[933] = 12'h00f;
rom[934] = 12'h000;
rom[935] = 12'h000;
rom[936] = 12'h000;
rom[937] = 12'h000;
rom[938] = 12'h007;
rom[939] = 12'h007;
rom[940] = 12'h000;
rom[941] = 12'h000;
rom[942] = 12'h007;
rom[943] = 12'h007;
rom[944] = 12'h000;
rom[945] = 12'h000;
rom[946] = 12'h000;
rom[947] = 12'h000;
rom[948] = 12'h000;
rom[949] = 12'h000;
rom[950] = 12'h000;
rom[951] = 12'h000;
rom[952] = 12'h000;
rom[953] = 12'h000;
rom[954] = 12'h00f;
rom[955] = 12'h00f;
rom[956] = 12'h00f;
rom[957] = 12'h00f;
rom[958] = 12'h00f;
rom[959] = 12'h00f;
rom[960] = 12'h000;
rom[961] = 12'h000;
rom[962] = 12'h000;
rom[963] = 12'h000;
rom[964] = 12'h007;
rom[965] = 12'h007;
rom[966] = 12'h000;
rom[967] = 12'h000;
rom[968] = 12'h007;
rom[969] = 12'h007;
rom[970] = 12'h000;
rom[971] = 12'h000;
rom[972] = 12'h000;
rom[973] = 12'h000;
rom[974] = 12'h000;
rom[975] = 12'h000;
rom[976] = 12'h000;
rom[977] = 12'h000;
rom[978] = 12'h000;
rom[979] = 12'h000;
rom[980] = 12'h00f;
rom[981] = 12'h00f;
rom[982] = 12'h00f;
rom[983] = 12'h00f;
rom[984] = 12'h00f;
rom[985] = 12'h00f;
rom[986] = 12'h000;
rom[987] = 12'h000;
rom[988] = 12'h000;
rom[989] = 12'h000;
rom[990] = 12'h000;
rom[991] = 12'h000;
rom[992] = 12'h007;
rom[993] = 12'h007;
rom[994] = 12'h000;
rom[995] = 12'h000;
rom[996] = 12'h00f;
rom[997] = 12'h00f;
rom[998] = 12'h00f;
rom[999] = 12'h00f;
rom[1000] = 12'h00f;
rom[1001] = 12'h00f;
rom[1002] = 12'h00f;
rom[1003] = 12'h00f;
rom[1004] = 12'h00f;
rom[1005] = 12'h00f;
rom[1006] = 12'h000;
rom[1007] = 12'h000;
rom[1008] = 12'h00f;
rom[1009] = 12'h00f;
rom[1010] = 12'h00f;
rom[1011] = 12'h00f;
rom[1012] = 12'h000;
rom[1013] = 12'h000;
rom[1014] = 12'h000;
rom[1015] = 12'h000;
rom[1016] = 12'h000;
rom[1017] = 12'h000;
rom[1018] = 12'h007;
rom[1019] = 12'h007;
rom[1020] = 12'h000;
rom[1021] = 12'h000;
rom[1022] = 12'h00f;
rom[1023] = 12'h00f;
rom[1024] = 12'h00f;
rom[1025] = 12'h00f;
rom[1026] = 12'h00f;
rom[1027] = 12'h00f;
rom[1028] = 12'h00f;
rom[1029] = 12'h00f;
rom[1030] = 12'h00f;
rom[1031] = 12'h00f;
rom[1032] = 12'h000;
rom[1033] = 12'h000;
rom[1034] = 12'h00f;
rom[1035] = 12'h00f;
rom[1036] = 12'h00f;
rom[1037] = 12'h00f;
rom[1038] = 12'h000;
rom[1039] = 12'h000;
rom[1040] = 12'h000;
rom[1041] = 12'h000;
rom[1042] = 12'h007;
rom[1043] = 12'h007;
rom[1044] = 12'h000;
rom[1045] = 12'h000;
rom[1046] = 12'h00f;
rom[1047] = 12'h00f;
rom[1048] = 12'h00f;
rom[1049] = 12'h00f;
rom[1050] = 12'h00f;
rom[1051] = 12'h00f;
rom[1052] = 12'h00f;
rom[1053] = 12'h00f;
rom[1054] = 12'h00f;
rom[1055] = 12'h00f;
rom[1056] = 12'h00f;
rom[1057] = 12'h00f;
rom[1058] = 12'h00f;
rom[1059] = 12'h00f;
rom[1060] = 12'h000;
rom[1061] = 12'h000;
rom[1062] = 12'h00f;
rom[1063] = 12'h00f;
rom[1064] = 12'h000;
rom[1065] = 12'h000;
rom[1066] = 12'h000;
rom[1067] = 12'h000;
rom[1068] = 12'h007;
rom[1069] = 12'h007;
rom[1070] = 12'h000;
rom[1071] = 12'h000;
rom[1072] = 12'h00f;
rom[1073] = 12'h00f;
rom[1074] = 12'h00f;
rom[1075] = 12'h00f;
rom[1076] = 12'h00f;
rom[1077] = 12'h00f;
rom[1078] = 12'h00f;
rom[1079] = 12'h00f;
rom[1080] = 12'h00f;
rom[1081] = 12'h00f;
rom[1082] = 12'h00f;
rom[1083] = 12'h00f;
rom[1084] = 12'h00f;
rom[1085] = 12'h00f;
rom[1086] = 12'h000;
rom[1087] = 12'h000;
rom[1088] = 12'h00f;
rom[1089] = 12'h00f;
rom[1090] = 12'h000;
rom[1091] = 12'h000;
rom[1092] = 12'h000;
rom[1093] = 12'h000;
rom[1094] = 12'h000;
rom[1095] = 12'h000;
rom[1096] = 12'h00f;
rom[1097] = 12'h00f;
rom[1098] = 12'h00f;
rom[1099] = 12'h00f;
rom[1100] = 12'h00f;
rom[1101] = 12'h00f;
rom[1102] = 12'h00f;
rom[1103] = 12'h00f;
rom[1104] = 12'h00f;
rom[1105] = 12'h00f;
rom[1106] = 12'h00f;
rom[1107] = 12'h00f;
rom[1108] = 12'h00f;
rom[1109] = 12'h00f;
rom[1110] = 12'h00f;
rom[1111] = 12'h00f;
rom[1112] = 12'h00f;
rom[1113] = 12'h00f;
rom[1114] = 12'h000;
rom[1115] = 12'h000;
rom[1116] = 12'h000;
rom[1117] = 12'h000;
rom[1118] = 12'h000;
rom[1119] = 12'h000;
rom[1120] = 12'h000;
rom[1121] = 12'h000;
rom[1122] = 12'h00f;
rom[1123] = 12'h00f;
rom[1124] = 12'h00f;
rom[1125] = 12'h00f;
rom[1126] = 12'h00f;
rom[1127] = 12'h00f;
rom[1128] = 12'h00f;
rom[1129] = 12'h00f;
rom[1130] = 12'h00f;
rom[1131] = 12'h00f;
rom[1132] = 12'h00f;
rom[1133] = 12'h00f;
rom[1134] = 12'h00f;
rom[1135] = 12'h00f;
rom[1136] = 12'h00f;
rom[1137] = 12'h00f;
rom[1138] = 12'h00f;
rom[1139] = 12'h00f;
rom[1140] = 12'h000;
rom[1141] = 12'h000;
rom[1142] = 12'h000;
rom[1143] = 12'h000;
rom[1144] = 12'h000;
rom[1145] = 12'h000;
rom[1146] = 12'h000;
rom[1147] = 12'h000;
rom[1148] = 12'h000;
rom[1149] = 12'h000;
rom[1150] = 12'h000;
rom[1151] = 12'h000;
rom[1152] = 12'h000;
rom[1153] = 12'h000;
rom[1154] = 12'h000;
rom[1155] = 12'h000;
rom[1156] = 12'h000;
rom[1157] = 12'h000;
rom[1158] = 12'h000;
rom[1159] = 12'h000;
rom[1160] = 12'h000;
rom[1161] = 12'h000;
rom[1162] = 12'h000;
rom[1163] = 12'h000;
rom[1164] = 12'h000;
rom[1165] = 12'h000;
rom[1166] = 12'h000;
rom[1167] = 12'h000;
rom[1168] = 12'h000;
rom[1169] = 12'h000;
rom[1170] = 12'h000;
rom[1171] = 12'h000;
rom[1172] = 12'h000;
rom[1173] = 12'h000;
rom[1174] = 12'h000;
rom[1175] = 12'h000;
rom[1176] = 12'h000;
rom[1177] = 12'h000;
rom[1178] = 12'h000;
rom[1179] = 12'h000;
rom[1180] = 12'h000;
rom[1181] = 12'h000;
rom[1182] = 12'h000;
rom[1183] = 12'h000;
rom[1184] = 12'h000;
rom[1185] = 12'h000;
rom[1186] = 12'h000;
rom[1187] = 12'h000;
rom[1188] = 12'h000;
rom[1189] = 12'h000;
rom[1190] = 12'h000;
rom[1191] = 12'h000;
rom[1192] = 12'h000;
rom[1193] = 12'h000;
rom[1194] = 12'h000;
rom[1195] = 12'h000;

  end
  endmodule

    module dash_rom (                       //шесть
  input  wire    [13:0]     addr,
  output wire    [11:0]     word
);

  logic [11:0] rom [(46 * 26)];

  assign word = rom[addr];

  initial begin
rom[0] = 12'h000;
rom[1] = 12'h000;
rom[2] = 12'h000;
rom[3] = 12'h000;
rom[4] = 12'h000;
rom[5] = 12'h000;
rom[6] = 12'h000;
rom[7] = 12'h000;
rom[8] = 12'h000;
rom[9] = 12'h000;
rom[10] = 12'h000;
rom[11] = 12'h000;
rom[12] = 12'h000;
rom[13] = 12'h000;
rom[14] = 12'h000;
rom[15] = 12'h000;
rom[16] = 12'h000;
rom[17] = 12'h000;
rom[18] = 12'h000;
rom[19] = 12'h000;
rom[20] = 12'h000;
rom[21] = 12'h000;
rom[22] = 12'h000;
rom[23] = 12'h000;
rom[24] = 12'h000;
rom[25] = 12'h000;
rom[26] = 12'h000;
rom[27] = 12'h000;
rom[28] = 12'h000;
rom[29] = 12'h000;
rom[30] = 12'h000;
rom[31] = 12'h000;
rom[32] = 12'h000;
rom[33] = 12'h000;
rom[34] = 12'h000;
rom[35] = 12'h000;
rom[36] = 12'h000;
rom[37] = 12'h000;
rom[38] = 12'h000;
rom[39] = 12'h000;
rom[40] = 12'h000;
rom[41] = 12'h000;
rom[42] = 12'h000;
rom[43] = 12'h000;
rom[44] = 12'h000;
rom[45] = 12'h000;
rom[46] = 12'h000;
rom[47] = 12'h000;
rom[48] = 12'h000;
rom[49] = 12'h000;
rom[50] = 12'h000;
rom[51] = 12'h000;
rom[52] = 12'h000;
rom[53] = 12'h000;
rom[54] = 12'h000;
rom[55] = 12'h000;
rom[56] = 12'h00f;
rom[57] = 12'h00f;
rom[58] = 12'h00f;
rom[59] = 12'h00f;
rom[60] = 12'h00f;
rom[61] = 12'h00f;
rom[62] = 12'h00f;
rom[63] = 12'h00f;
rom[64] = 12'h00f;
rom[65] = 12'h00f;
rom[66] = 12'h00f;
rom[67] = 12'h00f;
rom[68] = 12'h00f;
rom[69] = 12'h00f;
rom[70] = 12'h00f;
rom[71] = 12'h00f;
rom[72] = 12'h00f;
rom[73] = 12'h00f;
rom[74] = 12'h000;
rom[75] = 12'h000;
rom[76] = 12'h000;
rom[77] = 12'h000;
rom[78] = 12'h000;
rom[79] = 12'h000;
rom[80] = 12'h000;
rom[81] = 12'h000;
rom[82] = 12'h00f;
rom[83] = 12'h00f;
rom[84] = 12'h00f;
rom[85] = 12'h00f;
rom[86] = 12'h00f;
rom[87] = 12'h00f;
rom[88] = 12'h00f;
rom[89] = 12'h00f;
rom[90] = 12'h00f;
rom[91] = 12'h00f;
rom[92] = 12'h00f;
rom[93] = 12'h00f;
rom[94] = 12'h00f;
rom[95] = 12'h00f;
rom[96] = 12'h00f;
rom[97] = 12'h00f;
rom[98] = 12'h00f;
rom[99] = 12'h00f;
rom[100] = 12'h000;
rom[101] = 12'h000;
rom[102] = 12'h000;
rom[103] = 12'h000;
rom[104] = 12'h000;
rom[105] = 12'h000;
rom[106] = 12'h00f;
rom[107] = 12'h00f;
rom[108] = 12'h000;
rom[109] = 12'h000;
rom[110] = 12'h00f;
rom[111] = 12'h00f;
rom[112] = 12'h00f;
rom[113] = 12'h00f;
rom[114] = 12'h00f;
rom[115] = 12'h00f;
rom[116] = 12'h00f;
rom[117] = 12'h00f;
rom[118] = 12'h00f;
rom[119] = 12'h00f;
rom[120] = 12'h00f;
rom[121] = 12'h00f;
rom[122] = 12'h00f;
rom[123] = 12'h00f;
rom[124] = 12'h000;
rom[125] = 12'h000;
rom[126] = 12'h007;
rom[127] = 12'h007;
rom[128] = 12'h000;
rom[129] = 12'h000;
rom[130] = 12'h000;
rom[131] = 12'h000;
rom[132] = 12'h00f;
rom[133] = 12'h00f;
rom[134] = 12'h000;
rom[135] = 12'h000;
rom[136] = 12'h00f;
rom[137] = 12'h00f;
rom[138] = 12'h00f;
rom[139] = 12'h00f;
rom[140] = 12'h00f;
rom[141] = 12'h00f;
rom[142] = 12'h00f;
rom[143] = 12'h00f;
rom[144] = 12'h00f;
rom[145] = 12'h00f;
rom[146] = 12'h00f;
rom[147] = 12'h00f;
rom[148] = 12'h00f;
rom[149] = 12'h00f;
rom[150] = 12'h000;
rom[151] = 12'h000;
rom[152] = 12'h007;
rom[153] = 12'h007;
rom[154] = 12'h000;
rom[155] = 12'h000;
rom[156] = 12'h000;
rom[157] = 12'h000;
rom[158] = 12'h00f;
rom[159] = 12'h00f;
rom[160] = 12'h00f;
rom[161] = 12'h00f;
rom[162] = 12'h000;
rom[163] = 12'h000;
rom[164] = 12'h00f;
rom[165] = 12'h00f;
rom[166] = 12'h00f;
rom[167] = 12'h00f;
rom[168] = 12'h00f;
rom[169] = 12'h00f;
rom[170] = 12'h00f;
rom[171] = 12'h00f;
rom[172] = 12'h00f;
rom[173] = 12'h00f;
rom[174] = 12'h000;
rom[175] = 12'h000;
rom[176] = 12'h007;
rom[177] = 12'h007;
rom[178] = 12'h000;
rom[179] = 12'h000;
rom[180] = 12'h000;
rom[181] = 12'h000;
rom[182] = 12'h000;
rom[183] = 12'h000;
rom[184] = 12'h00f;
rom[185] = 12'h00f;
rom[186] = 12'h00f;
rom[187] = 12'h00f;
rom[188] = 12'h000;
rom[189] = 12'h000;
rom[190] = 12'h00f;
rom[191] = 12'h00f;
rom[192] = 12'h00f;
rom[193] = 12'h00f;
rom[194] = 12'h00f;
rom[195] = 12'h00f;
rom[196] = 12'h00f;
rom[197] = 12'h00f;
rom[198] = 12'h00f;
rom[199] = 12'h00f;
rom[200] = 12'h000;
rom[201] = 12'h000;
rom[202] = 12'h007;
rom[203] = 12'h007;
rom[204] = 12'h000;
rom[205] = 12'h000;
rom[206] = 12'h000;
rom[207] = 12'h000;
rom[208] = 12'h000;
rom[209] = 12'h000;
rom[210] = 12'h00f;
rom[211] = 12'h00f;
rom[212] = 12'h00f;
rom[213] = 12'h00f;
rom[214] = 12'h00f;
rom[215] = 12'h00f;
rom[216] = 12'h000;
rom[217] = 12'h000;
rom[218] = 12'h000;
rom[219] = 12'h000;
rom[220] = 12'h000;
rom[221] = 12'h000;
rom[222] = 12'h000;
rom[223] = 12'h000;
rom[224] = 12'h000;
rom[225] = 12'h000;
rom[226] = 12'h007;
rom[227] = 12'h007;
rom[228] = 12'h000;
rom[229] = 12'h000;
rom[230] = 12'h007;
rom[231] = 12'h007;
rom[232] = 12'h000;
rom[233] = 12'h000;
rom[234] = 12'h000;
rom[235] = 12'h000;
rom[236] = 12'h00f;
rom[237] = 12'h00f;
rom[238] = 12'h00f;
rom[239] = 12'h00f;
rom[240] = 12'h00f;
rom[241] = 12'h00f;
rom[242] = 12'h000;
rom[243] = 12'h000;
rom[244] = 12'h000;
rom[245] = 12'h000;
rom[246] = 12'h000;
rom[247] = 12'h000;
rom[248] = 12'h000;
rom[249] = 12'h000;
rom[250] = 12'h000;
rom[251] = 12'h000;
rom[252] = 12'h007;
rom[253] = 12'h007;
rom[254] = 12'h000;
rom[255] = 12'h000;
rom[256] = 12'h007;
rom[257] = 12'h007;
rom[258] = 12'h000;
rom[259] = 12'h000;
rom[260] = 12'h000;
rom[261] = 12'h000;
rom[262] = 12'h00f;
rom[263] = 12'h00f;
rom[264] = 12'h00f;
rom[265] = 12'h00f;
rom[266] = 12'h00f;
rom[267] = 12'h00f;
rom[268] = 12'h000;
rom[269] = 12'h000;
rom[270] = 12'h000;
rom[271] = 12'h000;
rom[272] = 12'h000;
rom[273] = 12'h000;
rom[274] = 12'h000;
rom[275] = 12'h000;
rom[276] = 12'h000;
rom[277] = 12'h000;
rom[278] = 12'h000;
rom[279] = 12'h000;
rom[280] = 12'h007;
rom[281] = 12'h007;
rom[282] = 12'h000;
rom[283] = 12'h000;
rom[284] = 12'h000;
rom[285] = 12'h000;
rom[286] = 12'h000;
rom[287] = 12'h000;
rom[288] = 12'h00f;
rom[289] = 12'h00f;
rom[290] = 12'h00f;
rom[291] = 12'h00f;
rom[292] = 12'h00f;
rom[293] = 12'h00f;
rom[294] = 12'h000;
rom[295] = 12'h000;
rom[296] = 12'h000;
rom[297] = 12'h000;
rom[298] = 12'h000;
rom[299] = 12'h000;
rom[300] = 12'h000;
rom[301] = 12'h000;
rom[302] = 12'h000;
rom[303] = 12'h000;
rom[304] = 12'h000;
rom[305] = 12'h000;
rom[306] = 12'h007;
rom[307] = 12'h007;
rom[308] = 12'h000;
rom[309] = 12'h000;
rom[310] = 12'h000;
rom[311] = 12'h000;
rom[312] = 12'h000;
rom[313] = 12'h000;
rom[314] = 12'h00f;
rom[315] = 12'h00f;
rom[316] = 12'h00f;
rom[317] = 12'h00f;
rom[318] = 12'h00f;
rom[319] = 12'h00f;
rom[320] = 12'h000;
rom[321] = 12'h000;
rom[322] = 12'h000;
rom[323] = 12'h000;
rom[324] = 12'h000;
rom[325] = 12'h000;
rom[326] = 12'h000;
rom[327] = 12'h000;
rom[328] = 12'h000;
rom[329] = 12'h000;
rom[330] = 12'h007;
rom[331] = 12'h007;
rom[332] = 12'h000;
rom[333] = 12'h000;
rom[334] = 12'h007;
rom[335] = 12'h007;
rom[336] = 12'h000;
rom[337] = 12'h000;
rom[338] = 12'h000;
rom[339] = 12'h000;
rom[340] = 12'h00f;
rom[341] = 12'h00f;
rom[342] = 12'h00f;
rom[343] = 12'h00f;
rom[344] = 12'h00f;
rom[345] = 12'h00f;
rom[346] = 12'h000;
rom[347] = 12'h000;
rom[348] = 12'h000;
rom[349] = 12'h000;
rom[350] = 12'h000;
rom[351] = 12'h000;
rom[352] = 12'h000;
rom[353] = 12'h000;
rom[354] = 12'h000;
rom[355] = 12'h000;
rom[356] = 12'h007;
rom[357] = 12'h007;
rom[358] = 12'h000;
rom[359] = 12'h000;
rom[360] = 12'h007;
rom[361] = 12'h007;
rom[362] = 12'h000;
rom[363] = 12'h000;
rom[364] = 12'h000;
rom[365] = 12'h000;
rom[366] = 12'h00f;
rom[367] = 12'h00f;
rom[368] = 12'h00f;
rom[369] = 12'h00f;
rom[370] = 12'h00f;
rom[371] = 12'h00f;
rom[372] = 12'h000;
rom[373] = 12'h000;
rom[374] = 12'h000;
rom[375] = 12'h000;
rom[376] = 12'h000;
rom[377] = 12'h000;
rom[378] = 12'h000;
rom[379] = 12'h000;
rom[380] = 12'h000;
rom[381] = 12'h000;
rom[382] = 12'h000;
rom[383] = 12'h000;
rom[384] = 12'h007;
rom[385] = 12'h007;
rom[386] = 12'h000;
rom[387] = 12'h000;
rom[388] = 12'h000;
rom[389] = 12'h000;
rom[390] = 12'h000;
rom[391] = 12'h000;
rom[392] = 12'h00f;
rom[393] = 12'h00f;
rom[394] = 12'h00f;
rom[395] = 12'h00f;
rom[396] = 12'h00f;
rom[397] = 12'h00f;
rom[398] = 12'h000;
rom[399] = 12'h000;
rom[400] = 12'h000;
rom[401] = 12'h000;
rom[402] = 12'h000;
rom[403] = 12'h000;
rom[404] = 12'h000;
rom[405] = 12'h000;
rom[406] = 12'h000;
rom[407] = 12'h000;
rom[408] = 12'h000;
rom[409] = 12'h000;
rom[410] = 12'h007;
rom[411] = 12'h007;
rom[412] = 12'h000;
rom[413] = 12'h000;
rom[414] = 12'h000;
rom[415] = 12'h000;
rom[416] = 12'h000;
rom[417] = 12'h000;
rom[418] = 12'h00f;
rom[419] = 12'h00f;
rom[420] = 12'h00f;
rom[421] = 12'h00f;
rom[422] = 12'h00f;
rom[423] = 12'h00f;
rom[424] = 12'h000;
rom[425] = 12'h000;
rom[426] = 12'h000;
rom[427] = 12'h000;
rom[428] = 12'h000;
rom[429] = 12'h000;
rom[430] = 12'h000;
rom[431] = 12'h000;
rom[432] = 12'h000;
rom[433] = 12'h000;
rom[434] = 12'h007;
rom[435] = 12'h007;
rom[436] = 12'h000;
rom[437] = 12'h000;
rom[438] = 12'h007;
rom[439] = 12'h007;
rom[440] = 12'h000;
rom[441] = 12'h000;
rom[442] = 12'h000;
rom[443] = 12'h000;
rom[444] = 12'h00f;
rom[445] = 12'h00f;
rom[446] = 12'h00f;
rom[447] = 12'h00f;
rom[448] = 12'h00f;
rom[449] = 12'h00f;
rom[450] = 12'h000;
rom[451] = 12'h000;
rom[452] = 12'h000;
rom[453] = 12'h000;
rom[454] = 12'h000;
rom[455] = 12'h000;
rom[456] = 12'h000;
rom[457] = 12'h000;
rom[458] = 12'h000;
rom[459] = 12'h000;
rom[460] = 12'h007;
rom[461] = 12'h007;
rom[462] = 12'h000;
rom[463] = 12'h000;
rom[464] = 12'h007;
rom[465] = 12'h007;
rom[466] = 12'h000;
rom[467] = 12'h000;
rom[468] = 12'h000;
rom[469] = 12'h000;
rom[470] = 12'h00f;
rom[471] = 12'h00f;
rom[472] = 12'h00f;
rom[473] = 12'h00f;
rom[474] = 12'h000;
rom[475] = 12'h000;
rom[476] = 12'h000;
rom[477] = 12'h000;
rom[478] = 12'h000;
rom[479] = 12'h000;
rom[480] = 12'h000;
rom[481] = 12'h000;
rom[482] = 12'h000;
rom[483] = 12'h000;
rom[484] = 12'h000;
rom[485] = 12'h000;
rom[486] = 12'h000;
rom[487] = 12'h000;
rom[488] = 12'h007;
rom[489] = 12'h007;
rom[490] = 12'h000;
rom[491] = 12'h000;
rom[492] = 12'h000;
rom[493] = 12'h000;
rom[494] = 12'h000;
rom[495] = 12'h000;
rom[496] = 12'h00f;
rom[497] = 12'h00f;
rom[498] = 12'h00f;
rom[499] = 12'h00f;
rom[500] = 12'h000;
rom[501] = 12'h000;
rom[502] = 12'h000;
rom[503] = 12'h000;
rom[504] = 12'h000;
rom[505] = 12'h000;
rom[506] = 12'h000;
rom[507] = 12'h000;
rom[508] = 12'h000;
rom[509] = 12'h000;
rom[510] = 12'h000;
rom[511] = 12'h000;
rom[512] = 12'h000;
rom[513] = 12'h000;
rom[514] = 12'h007;
rom[515] = 12'h007;
rom[516] = 12'h000;
rom[517] = 12'h000;
rom[518] = 12'h000;
rom[519] = 12'h000;
rom[520] = 12'h000;
rom[521] = 12'h000;
rom[522] = 12'h00f;
rom[523] = 12'h00f;
rom[524] = 12'h000;
rom[525] = 12'h000;
rom[526] = 12'h00f;
rom[527] = 12'h00f;
rom[528] = 12'h00f;
rom[529] = 12'h00f;
rom[530] = 12'h00f;
rom[531] = 12'h00f;
rom[532] = 12'h00f;
rom[533] = 12'h00f;
rom[534] = 12'h00f;
rom[535] = 12'h00f;
rom[536] = 12'h00f;
rom[537] = 12'h00f;
rom[538] = 12'h00f;
rom[539] = 12'h00f;
rom[540] = 12'h000;
rom[541] = 12'h000;
rom[542] = 12'h007;
rom[543] = 12'h007;
rom[544] = 12'h000;
rom[545] = 12'h000;
rom[546] = 12'h000;
rom[547] = 12'h000;
rom[548] = 12'h00f;
rom[549] = 12'h00f;
rom[550] = 12'h000;
rom[551] = 12'h000;
rom[552] = 12'h00f;
rom[553] = 12'h00f;
rom[554] = 12'h00f;
rom[555] = 12'h00f;
rom[556] = 12'h00f;
rom[557] = 12'h00f;
rom[558] = 12'h00f;
rom[559] = 12'h00f;
rom[560] = 12'h00f;
rom[561] = 12'h00f;
rom[562] = 12'h00f;
rom[563] = 12'h00f;
rom[564] = 12'h00f;
rom[565] = 12'h00f;
rom[566] = 12'h000;
rom[567] = 12'h000;
rom[568] = 12'h007;
rom[569] = 12'h007;
rom[570] = 12'h000;
rom[571] = 12'h000;
rom[572] = 12'h000;
rom[573] = 12'h000;
rom[574] = 12'h000;
rom[575] = 12'h000;
rom[576] = 12'h00f;
rom[577] = 12'h00f;
rom[578] = 12'h00f;
rom[579] = 12'h00f;
rom[580] = 12'h00f;
rom[581] = 12'h00f;
rom[582] = 12'h00f;
rom[583] = 12'h00f;
rom[584] = 12'h00f;
rom[585] = 12'h00f;
rom[586] = 12'h00f;
rom[587] = 12'h00f;
rom[588] = 12'h00f;
rom[589] = 12'h00f;
rom[590] = 12'h00f;
rom[591] = 12'h00f;
rom[592] = 12'h00f;
rom[593] = 12'h00f;
rom[594] = 12'h000;
rom[595] = 12'h000;
rom[596] = 12'h000;
rom[597] = 12'h000;
rom[598] = 12'h000;
rom[599] = 12'h000;
rom[600] = 12'h000;
rom[601] = 12'h000;
rom[602] = 12'h00f;
rom[603] = 12'h00f;
rom[604] = 12'h00f;
rom[605] = 12'h00f;
rom[606] = 12'h00f;
rom[607] = 12'h00f;
rom[608] = 12'h00f;
rom[609] = 12'h00f;
rom[610] = 12'h00f;
rom[611] = 12'h00f;
rom[612] = 12'h00f;
rom[613] = 12'h00f;
rom[614] = 12'h00f;
rom[615] = 12'h00f;
rom[616] = 12'h00f;
rom[617] = 12'h00f;
rom[618] = 12'h00f;
rom[619] = 12'h00f;
rom[620] = 12'h000;
rom[621] = 12'h000;
rom[622] = 12'h000;
rom[623] = 12'h000;
rom[624] = 12'h000;
rom[625] = 12'h000;
rom[626] = 12'h00f;
rom[627] = 12'h00f;
rom[628] = 12'h000;
rom[629] = 12'h000;
rom[630] = 12'h00f;
rom[631] = 12'h00f;
rom[632] = 12'h00f;
rom[633] = 12'h00f;
rom[634] = 12'h00f;
rom[635] = 12'h00f;
rom[636] = 12'h00f;
rom[637] = 12'h00f;
rom[638] = 12'h00f;
rom[639] = 12'h00f;
rom[640] = 12'h00f;
rom[641] = 12'h00f;
rom[642] = 12'h00f;
rom[643] = 12'h00f;
rom[644] = 12'h000;
rom[645] = 12'h000;
rom[646] = 12'h00f;
rom[647] = 12'h00f;
rom[648] = 12'h000;
rom[649] = 12'h000;
rom[650] = 12'h000;
rom[651] = 12'h000;
rom[652] = 12'h00f;
rom[653] = 12'h00f;
rom[654] = 12'h000;
rom[655] = 12'h000;
rom[656] = 12'h00f;
rom[657] = 12'h00f;
rom[658] = 12'h00f;
rom[659] = 12'h00f;
rom[660] = 12'h00f;
rom[661] = 12'h00f;
rom[662] = 12'h00f;
rom[663] = 12'h00f;
rom[664] = 12'h00f;
rom[665] = 12'h00f;
rom[666] = 12'h00f;
rom[667] = 12'h00f;
rom[668] = 12'h00f;
rom[669] = 12'h00f;
rom[670] = 12'h000;
rom[671] = 12'h000;
rom[672] = 12'h00f;
rom[673] = 12'h00f;
rom[674] = 12'h000;
rom[675] = 12'h000;
rom[676] = 12'h000;
rom[677] = 12'h000;
rom[678] = 12'h00f;
rom[679] = 12'h00f;
rom[680] = 12'h00f;
rom[681] = 12'h00f;
rom[682] = 12'h000;
rom[683] = 12'h000;
rom[684] = 12'h000;
rom[685] = 12'h000;
rom[686] = 12'h000;
rom[687] = 12'h000;
rom[688] = 12'h000;
rom[689] = 12'h000;
rom[690] = 12'h000;
rom[691] = 12'h000;
rom[692] = 12'h000;
rom[693] = 12'h000;
rom[694] = 12'h000;
rom[695] = 12'h000;
rom[696] = 12'h00f;
rom[697] = 12'h00f;
rom[698] = 12'h00f;
rom[699] = 12'h00f;
rom[700] = 12'h000;
rom[701] = 12'h000;
rom[702] = 12'h000;
rom[703] = 12'h000;
rom[704] = 12'h00f;
rom[705] = 12'h00f;
rom[706] = 12'h00f;
rom[707] = 12'h00f;
rom[708] = 12'h000;
rom[709] = 12'h000;
rom[710] = 12'h000;
rom[711] = 12'h000;
rom[712] = 12'h000;
rom[713] = 12'h000;
rom[714] = 12'h000;
rom[715] = 12'h000;
rom[716] = 12'h000;
rom[717] = 12'h000;
rom[718] = 12'h000;
rom[719] = 12'h000;
rom[720] = 12'h000;
rom[721] = 12'h000;
rom[722] = 12'h00f;
rom[723] = 12'h00f;
rom[724] = 12'h00f;
rom[725] = 12'h00f;
rom[726] = 12'h000;
rom[727] = 12'h000;
rom[728] = 12'h000;
rom[729] = 12'h000;
rom[730] = 12'h00f;
rom[731] = 12'h00f;
rom[732] = 12'h00f;
rom[733] = 12'h00f;
rom[734] = 12'h00f;
rom[735] = 12'h00f;
rom[736] = 12'h000;
rom[737] = 12'h000;
rom[738] = 12'h000;
rom[739] = 12'h000;
rom[740] = 12'h000;
rom[741] = 12'h000;
rom[742] = 12'h000;
rom[743] = 12'h000;
rom[744] = 12'h000;
rom[745] = 12'h000;
rom[746] = 12'h00f;
rom[747] = 12'h00f;
rom[748] = 12'h00f;
rom[749] = 12'h00f;
rom[750] = 12'h00f;
rom[751] = 12'h00f;
rom[752] = 12'h000;
rom[753] = 12'h000;
rom[754] = 12'h000;
rom[755] = 12'h000;
rom[756] = 12'h00f;
rom[757] = 12'h00f;
rom[758] = 12'h00f;
rom[759] = 12'h00f;
rom[760] = 12'h00f;
rom[761] = 12'h00f;
rom[762] = 12'h000;
rom[763] = 12'h000;
rom[764] = 12'h000;
rom[765] = 12'h000;
rom[766] = 12'h000;
rom[767] = 12'h000;
rom[768] = 12'h000;
rom[769] = 12'h000;
rom[770] = 12'h000;
rom[771] = 12'h000;
rom[772] = 12'h00f;
rom[773] = 12'h00f;
rom[774] = 12'h00f;
rom[775] = 12'h00f;
rom[776] = 12'h00f;
rom[777] = 12'h00f;
rom[778] = 12'h000;
rom[779] = 12'h000;
rom[780] = 12'h000;
rom[781] = 12'h000;
rom[782] = 12'h00f;
rom[783] = 12'h00f;
rom[784] = 12'h00f;
rom[785] = 12'h00f;
rom[786] = 12'h00f;
rom[787] = 12'h00f;
rom[788] = 12'h000;
rom[789] = 12'h000;
rom[790] = 12'h000;
rom[791] = 12'h000;
rom[792] = 12'h000;
rom[793] = 12'h000;
rom[794] = 12'h000;
rom[795] = 12'h000;
rom[796] = 12'h000;
rom[797] = 12'h000;
rom[798] = 12'h00f;
rom[799] = 12'h00f;
rom[800] = 12'h00f;
rom[801] = 12'h00f;
rom[802] = 12'h00f;
rom[803] = 12'h00f;
rom[804] = 12'h000;
rom[805] = 12'h000;
rom[806] = 12'h000;
rom[807] = 12'h000;
rom[808] = 12'h00f;
rom[809] = 12'h00f;
rom[810] = 12'h00f;
rom[811] = 12'h00f;
rom[812] = 12'h00f;
rom[813] = 12'h00f;
rom[814] = 12'h000;
rom[815] = 12'h000;
rom[816] = 12'h000;
rom[817] = 12'h000;
rom[818] = 12'h000;
rom[819] = 12'h000;
rom[820] = 12'h000;
rom[821] = 12'h000;
rom[822] = 12'h000;
rom[823] = 12'h000;
rom[824] = 12'h00f;
rom[825] = 12'h00f;
rom[826] = 12'h00f;
rom[827] = 12'h00f;
rom[828] = 12'h00f;
rom[829] = 12'h00f;
rom[830] = 12'h000;
rom[831] = 12'h000;
rom[832] = 12'h000;
rom[833] = 12'h000;
rom[834] = 12'h00f;
rom[835] = 12'h00f;
rom[836] = 12'h00f;
rom[837] = 12'h00f;
rom[838] = 12'h00f;
rom[839] = 12'h00f;
rom[840] = 12'h000;
rom[841] = 12'h000;
rom[842] = 12'h000;
rom[843] = 12'h000;
rom[844] = 12'h000;
rom[845] = 12'h000;
rom[846] = 12'h000;
rom[847] = 12'h000;
rom[848] = 12'h000;
rom[849] = 12'h000;
rom[850] = 12'h00f;
rom[851] = 12'h00f;
rom[852] = 12'h00f;
rom[853] = 12'h00f;
rom[854] = 12'h00f;
rom[855] = 12'h00f;
rom[856] = 12'h000;
rom[857] = 12'h000;
rom[858] = 12'h000;
rom[859] = 12'h000;
rom[860] = 12'h00f;
rom[861] = 12'h00f;
rom[862] = 12'h00f;
rom[863] = 12'h00f;
rom[864] = 12'h00f;
rom[865] = 12'h00f;
rom[866] = 12'h000;
rom[867] = 12'h000;
rom[868] = 12'h000;
rom[869] = 12'h000;
rom[870] = 12'h000;
rom[871] = 12'h000;
rom[872] = 12'h000;
rom[873] = 12'h000;
rom[874] = 12'h000;
rom[875] = 12'h000;
rom[876] = 12'h00f;
rom[877] = 12'h00f;
rom[878] = 12'h00f;
rom[879] = 12'h00f;
rom[880] = 12'h00f;
rom[881] = 12'h00f;
rom[882] = 12'h000;
rom[883] = 12'h000;
rom[884] = 12'h000;
rom[885] = 12'h000;
rom[886] = 12'h00f;
rom[887] = 12'h00f;
rom[888] = 12'h00f;
rom[889] = 12'h00f;
rom[890] = 12'h00f;
rom[891] = 12'h00f;
rom[892] = 12'h000;
rom[893] = 12'h000;
rom[894] = 12'h000;
rom[895] = 12'h000;
rom[896] = 12'h000;
rom[897] = 12'h000;
rom[898] = 12'h000;
rom[899] = 12'h000;
rom[900] = 12'h000;
rom[901] = 12'h000;
rom[902] = 12'h00f;
rom[903] = 12'h00f;
rom[904] = 12'h00f;
rom[905] = 12'h00f;
rom[906] = 12'h00f;
rom[907] = 12'h00f;
rom[908] = 12'h000;
rom[909] = 12'h000;
rom[910] = 12'h000;
rom[911] = 12'h000;
rom[912] = 12'h00f;
rom[913] = 12'h00f;
rom[914] = 12'h00f;
rom[915] = 12'h00f;
rom[916] = 12'h00f;
rom[917] = 12'h00f;
rom[918] = 12'h000;
rom[919] = 12'h000;
rom[920] = 12'h000;
rom[921] = 12'h000;
rom[922] = 12'h000;
rom[923] = 12'h000;
rom[924] = 12'h000;
rom[925] = 12'h000;
rom[926] = 12'h000;
rom[927] = 12'h000;
rom[928] = 12'h00f;
rom[929] = 12'h00f;
rom[930] = 12'h00f;
rom[931] = 12'h00f;
rom[932] = 12'h00f;
rom[933] = 12'h00f;
rom[934] = 12'h000;
rom[935] = 12'h000;
rom[936] = 12'h000;
rom[937] = 12'h000;
rom[938] = 12'h00f;
rom[939] = 12'h00f;
rom[940] = 12'h00f;
rom[941] = 12'h00f;
rom[942] = 12'h00f;
rom[943] = 12'h00f;
rom[944] = 12'h000;
rom[945] = 12'h000;
rom[946] = 12'h000;
rom[947] = 12'h000;
rom[948] = 12'h000;
rom[949] = 12'h000;
rom[950] = 12'h000;
rom[951] = 12'h000;
rom[952] = 12'h000;
rom[953] = 12'h000;
rom[954] = 12'h00f;
rom[955] = 12'h00f;
rom[956] = 12'h00f;
rom[957] = 12'h00f;
rom[958] = 12'h00f;
rom[959] = 12'h00f;
rom[960] = 12'h000;
rom[961] = 12'h000;
rom[962] = 12'h000;
rom[963] = 12'h000;
rom[964] = 12'h00f;
rom[965] = 12'h00f;
rom[966] = 12'h00f;
rom[967] = 12'h00f;
rom[968] = 12'h00f;
rom[969] = 12'h00f;
rom[970] = 12'h000;
rom[971] = 12'h000;
rom[972] = 12'h000;
rom[973] = 12'h000;
rom[974] = 12'h000;
rom[975] = 12'h000;
rom[976] = 12'h000;
rom[977] = 12'h000;
rom[978] = 12'h000;
rom[979] = 12'h000;
rom[980] = 12'h00f;
rom[981] = 12'h00f;
rom[982] = 12'h00f;
rom[983] = 12'h00f;
rom[984] = 12'h00f;
rom[985] = 12'h00f;
rom[986] = 12'h000;
rom[987] = 12'h000;
rom[988] = 12'h000;
rom[989] = 12'h000;
rom[990] = 12'h00f;
rom[991] = 12'h00f;
rom[992] = 12'h00f;
rom[993] = 12'h00f;
rom[994] = 12'h000;
rom[995] = 12'h000;
rom[996] = 12'h00f;
rom[997] = 12'h00f;
rom[998] = 12'h00f;
rom[999] = 12'h00f;
rom[1000] = 12'h00f;
rom[1001] = 12'h00f;
rom[1002] = 12'h00f;
rom[1003] = 12'h00f;
rom[1004] = 12'h00f;
rom[1005] = 12'h00f;
rom[1006] = 12'h000;
rom[1007] = 12'h000;
rom[1008] = 12'h00f;
rom[1009] = 12'h00f;
rom[1010] = 12'h00f;
rom[1011] = 12'h00f;
rom[1012] = 12'h000;
rom[1013] = 12'h000;
rom[1014] = 12'h000;
rom[1015] = 12'h000;
rom[1016] = 12'h00f;
rom[1017] = 12'h00f;
rom[1018] = 12'h00f;
rom[1019] = 12'h00f;
rom[1020] = 12'h000;
rom[1021] = 12'h000;
rom[1022] = 12'h00f;
rom[1023] = 12'h00f;
rom[1024] = 12'h00f;
rom[1025] = 12'h00f;
rom[1026] = 12'h00f;
rom[1027] = 12'h00f;
rom[1028] = 12'h00f;
rom[1029] = 12'h00f;
rom[1030] = 12'h00f;
rom[1031] = 12'h00f;
rom[1032] = 12'h000;
rom[1033] = 12'h000;
rom[1034] = 12'h00f;
rom[1035] = 12'h00f;
rom[1036] = 12'h00f;
rom[1037] = 12'h00f;
rom[1038] = 12'h000;
rom[1039] = 12'h000;
rom[1040] = 12'h000;
rom[1041] = 12'h000;
rom[1042] = 12'h00f;
rom[1043] = 12'h00f;
rom[1044] = 12'h000;
rom[1045] = 12'h000;
rom[1046] = 12'h00f;
rom[1047] = 12'h00f;
rom[1048] = 12'h00f;
rom[1049] = 12'h00f;
rom[1050] = 12'h00f;
rom[1051] = 12'h00f;
rom[1052] = 12'h00f;
rom[1053] = 12'h00f;
rom[1054] = 12'h00f;
rom[1055] = 12'h00f;
rom[1056] = 12'h00f;
rom[1057] = 12'h00f;
rom[1058] = 12'h00f;
rom[1059] = 12'h00f;
rom[1060] = 12'h000;
rom[1061] = 12'h000;
rom[1062] = 12'h00f;
rom[1063] = 12'h00f;
rom[1064] = 12'h000;
rom[1065] = 12'h000;
rom[1066] = 12'h000;
rom[1067] = 12'h000;
rom[1068] = 12'h00f;
rom[1069] = 12'h00f;
rom[1070] = 12'h000;
rom[1071] = 12'h000;
rom[1072] = 12'h00f;
rom[1073] = 12'h00f;
rom[1074] = 12'h00f;
rom[1075] = 12'h00f;
rom[1076] = 12'h00f;
rom[1077] = 12'h00f;
rom[1078] = 12'h00f;
rom[1079] = 12'h00f;
rom[1080] = 12'h00f;
rom[1081] = 12'h00f;
rom[1082] = 12'h00f;
rom[1083] = 12'h00f;
rom[1084] = 12'h00f;
rom[1085] = 12'h00f;
rom[1086] = 12'h000;
rom[1087] = 12'h000;
rom[1088] = 12'h00f;
rom[1089] = 12'h00f;
rom[1090] = 12'h000;
rom[1091] = 12'h000;
rom[1092] = 12'h000;
rom[1093] = 12'h000;
rom[1094] = 12'h000;
rom[1095] = 12'h000;
rom[1096] = 12'h00f;
rom[1097] = 12'h00f;
rom[1098] = 12'h00f;
rom[1099] = 12'h00f;
rom[1100] = 12'h00f;
rom[1101] = 12'h00f;
rom[1102] = 12'h00f;
rom[1103] = 12'h00f;
rom[1104] = 12'h00f;
rom[1105] = 12'h00f;
rom[1106] = 12'h00f;
rom[1107] = 12'h00f;
rom[1108] = 12'h00f;
rom[1109] = 12'h00f;
rom[1110] = 12'h00f;
rom[1111] = 12'h00f;
rom[1112] = 12'h00f;
rom[1113] = 12'h00f;
rom[1114] = 12'h000;
rom[1115] = 12'h000;
rom[1116] = 12'h000;
rom[1117] = 12'h000;
rom[1118] = 12'h000;
rom[1119] = 12'h000;
rom[1120] = 12'h000;
rom[1121] = 12'h000;
rom[1122] = 12'h00f;
rom[1123] = 12'h00f;
rom[1124] = 12'h00f;
rom[1125] = 12'h00f;
rom[1126] = 12'h00f;
rom[1127] = 12'h00f;
rom[1128] = 12'h00f;
rom[1129] = 12'h00f;
rom[1130] = 12'h00f;
rom[1131] = 12'h00f;
rom[1132] = 12'h00f;
rom[1133] = 12'h00f;
rom[1134] = 12'h00f;
rom[1135] = 12'h00f;
rom[1136] = 12'h00f;
rom[1137] = 12'h00f;
rom[1138] = 12'h00f;
rom[1139] = 12'h00f;
rom[1140] = 12'h000;
rom[1141] = 12'h000;
rom[1142] = 12'h000;
rom[1143] = 12'h000;
rom[1144] = 12'h000;
rom[1145] = 12'h000;
rom[1146] = 12'h000;
rom[1147] = 12'h000;
rom[1148] = 12'h000;
rom[1149] = 12'h000;
rom[1150] = 12'h000;
rom[1151] = 12'h000;
rom[1152] = 12'h000;
rom[1153] = 12'h000;
rom[1154] = 12'h000;
rom[1155] = 12'h000;
rom[1156] = 12'h000;
rom[1157] = 12'h000;
rom[1158] = 12'h000;
rom[1159] = 12'h000;
rom[1160] = 12'h000;
rom[1161] = 12'h000;
rom[1162] = 12'h000;
rom[1163] = 12'h000;
rom[1164] = 12'h000;
rom[1165] = 12'h000;
rom[1166] = 12'h000;
rom[1167] = 12'h000;
rom[1168] = 12'h000;
rom[1169] = 12'h000;
rom[1170] = 12'h000;
rom[1171] = 12'h000;
rom[1172] = 12'h000;
rom[1173] = 12'h000;
rom[1174] = 12'h000;
rom[1175] = 12'h000;
rom[1176] = 12'h000;
rom[1177] = 12'h000;
rom[1178] = 12'h000;
rom[1179] = 12'h000;
rom[1180] = 12'h000;
rom[1181] = 12'h000;
rom[1182] = 12'h000;
rom[1183] = 12'h000;
rom[1184] = 12'h000;
rom[1185] = 12'h000;
rom[1186] = 12'h000;
rom[1187] = 12'h000;
rom[1188] = 12'h000;
rom[1189] = 12'h000;
rom[1190] = 12'h000;
rom[1191] = 12'h000;
rom[1192] = 12'h000;
rom[1193] = 12'h000;
rom[1194] = 12'h000;
rom[1195] = 12'h000;

  end
  endmodule

    module dash_rom (                       //семь
  input  wire    [13:0]     addr,
  output wire    [11:0]     word
);

  logic [11:0] rom [(46 * 26)];

  assign word = rom[addr];

  initial begin
rom[0] = 12'h000;
rom[1] = 12'h000;
rom[2] = 12'h000;
rom[3] = 12'h000;
rom[4] = 12'h000;
rom[5] = 12'h000;
rom[6] = 12'h000;
rom[7] = 12'h000;
rom[8] = 12'h000;
rom[9] = 12'h000;
rom[10] = 12'h000;
rom[11] = 12'h000;
rom[12] = 12'h000;
rom[13] = 12'h000;
rom[14] = 12'h000;
rom[15] = 12'h000;
rom[16] = 12'h000;
rom[17] = 12'h000;
rom[18] = 12'h000;
rom[19] = 12'h000;
rom[20] = 12'h000;
rom[21] = 12'h000;
rom[22] = 12'h000;
rom[23] = 12'h000;
rom[24] = 12'h000;
rom[25] = 12'h000;
rom[26] = 12'h000;
rom[27] = 12'h000;
rom[28] = 12'h000;
rom[29] = 12'h000;
rom[30] = 12'h000;
rom[31] = 12'h000;
rom[32] = 12'h000;
rom[33] = 12'h000;
rom[34] = 12'h000;
rom[35] = 12'h000;
rom[36] = 12'h000;
rom[37] = 12'h000;
rom[38] = 12'h000;
rom[39] = 12'h000;
rom[40] = 12'h000;
rom[41] = 12'h000;
rom[42] = 12'h000;
rom[43] = 12'h000;
rom[44] = 12'h000;
rom[45] = 12'h000;
rom[46] = 12'h000;
rom[47] = 12'h000;
rom[48] = 12'h000;
rom[49] = 12'h000;
rom[50] = 12'h000;
rom[51] = 12'h000;
rom[52] = 12'h000;
rom[53] = 12'h000;
rom[54] = 12'h000;
rom[55] = 12'h000;
rom[56] = 12'h00f;
rom[57] = 12'h00f;
rom[58] = 12'h00f;
rom[59] = 12'h00f;
rom[60] = 12'h00f;
rom[61] = 12'h00f;
rom[62] = 12'h00f;
rom[63] = 12'h00f;
rom[64] = 12'h00f;
rom[65] = 12'h00f;
rom[66] = 12'h00f;
rom[67] = 12'h00f;
rom[68] = 12'h00f;
rom[69] = 12'h00f;
rom[70] = 12'h00f;
rom[71] = 12'h00f;
rom[72] = 12'h00f;
rom[73] = 12'h00f;
rom[74] = 12'h000;
rom[75] = 12'h000;
rom[76] = 12'h000;
rom[77] = 12'h000;
rom[78] = 12'h000;
rom[79] = 12'h000;
rom[80] = 12'h000;
rom[81] = 12'h000;
rom[82] = 12'h00f;
rom[83] = 12'h00f;
rom[84] = 12'h00f;
rom[85] = 12'h00f;
rom[86] = 12'h00f;
rom[87] = 12'h00f;
rom[88] = 12'h00f;
rom[89] = 12'h00f;
rom[90] = 12'h00f;
rom[91] = 12'h00f;
rom[92] = 12'h00f;
rom[93] = 12'h00f;
rom[94] = 12'h00f;
rom[95] = 12'h00f;
rom[96] = 12'h00f;
rom[97] = 12'h00f;
rom[98] = 12'h00f;
rom[99] = 12'h00f;
rom[100] = 12'h000;
rom[101] = 12'h000;
rom[102] = 12'h000;
rom[103] = 12'h000;
rom[104] = 12'h000;
rom[105] = 12'h000;
rom[106] = 12'h007;
rom[107] = 12'h007;
rom[108] = 12'h000;
rom[109] = 12'h000;
rom[110] = 12'h00f;
rom[111] = 12'h00f;
rom[112] = 12'h00f;
rom[113] = 12'h00f;
rom[114] = 12'h00f;
rom[115] = 12'h00f;
rom[116] = 12'h00f;
rom[117] = 12'h00f;
rom[118] = 12'h00f;
rom[119] = 12'h00f;
rom[120] = 12'h00f;
rom[121] = 12'h00f;
rom[122] = 12'h00f;
rom[123] = 12'h00f;
rom[124] = 12'h000;
rom[125] = 12'h000;
rom[126] = 12'h00f;
rom[127] = 12'h00f;
rom[128] = 12'h000;
rom[129] = 12'h000;
rom[130] = 12'h000;
rom[131] = 12'h000;
rom[132] = 12'h007;
rom[133] = 12'h007;
rom[134] = 12'h000;
rom[135] = 12'h000;
rom[136] = 12'h00f;
rom[137] = 12'h00f;
rom[138] = 12'h00f;
rom[139] = 12'h00f;
rom[140] = 12'h00f;
rom[141] = 12'h00f;
rom[142] = 12'h00f;
rom[143] = 12'h00f;
rom[144] = 12'h00f;
rom[145] = 12'h00f;
rom[146] = 12'h00f;
rom[147] = 12'h00f;
rom[148] = 12'h00f;
rom[149] = 12'h00f;
rom[150] = 12'h000;
rom[151] = 12'h000;
rom[152] = 12'h00f;
rom[153] = 12'h00f;
rom[154] = 12'h000;
rom[155] = 12'h000;
rom[156] = 12'h000;
rom[157] = 12'h000;
rom[158] = 12'h000;
rom[159] = 12'h000;
rom[160] = 12'h007;
rom[161] = 12'h007;
rom[162] = 12'h000;
rom[163] = 12'h000;
rom[164] = 12'h00f;
rom[165] = 12'h00f;
rom[166] = 12'h00f;
rom[167] = 12'h00f;
rom[168] = 12'h00f;
rom[169] = 12'h00f;
rom[170] = 12'h00f;
rom[171] = 12'h00f;
rom[172] = 12'h00f;
rom[173] = 12'h00f;
rom[174] = 12'h000;
rom[175] = 12'h000;
rom[176] = 12'h00f;
rom[177] = 12'h00f;
rom[178] = 12'h00f;
rom[179] = 12'h00f;
rom[180] = 12'h000;
rom[181] = 12'h000;
rom[182] = 12'h000;
rom[183] = 12'h000;
rom[184] = 12'h000;
rom[185] = 12'h000;
rom[186] = 12'h007;
rom[187] = 12'h007;
rom[188] = 12'h000;
rom[189] = 12'h000;
rom[190] = 12'h00f;
rom[191] = 12'h00f;
rom[192] = 12'h00f;
rom[193] = 12'h00f;
rom[194] = 12'h00f;
rom[195] = 12'h00f;
rom[196] = 12'h00f;
rom[197] = 12'h00f;
rom[198] = 12'h00f;
rom[199] = 12'h00f;
rom[200] = 12'h000;
rom[201] = 12'h000;
rom[202] = 12'h00f;
rom[203] = 12'h00f;
rom[204] = 12'h00f;
rom[205] = 12'h00f;
rom[206] = 12'h000;
rom[207] = 12'h000;
rom[208] = 12'h000;
rom[209] = 12'h000;
rom[210] = 12'h007;
rom[211] = 12'h007;
rom[212] = 12'h000;
rom[213] = 12'h000;
rom[214] = 12'h007;
rom[215] = 12'h007;
rom[216] = 12'h000;
rom[217] = 12'h000;
rom[218] = 12'h000;
rom[219] = 12'h000;
rom[220] = 12'h000;
rom[221] = 12'h000;
rom[222] = 12'h000;
rom[223] = 12'h000;
rom[224] = 12'h000;
rom[225] = 12'h000;
rom[226] = 12'h00f;
rom[227] = 12'h00f;
rom[228] = 12'h00f;
rom[229] = 12'h00f;
rom[230] = 12'h00f;
rom[231] = 12'h00f;
rom[232] = 12'h000;
rom[233] = 12'h000;
rom[234] = 12'h000;
rom[235] = 12'h000;
rom[236] = 12'h007;
rom[237] = 12'h007;
rom[238] = 12'h000;
rom[239] = 12'h000;
rom[240] = 12'h007;
rom[241] = 12'h007;
rom[242] = 12'h000;
rom[243] = 12'h000;
rom[244] = 12'h000;
rom[245] = 12'h000;
rom[246] = 12'h000;
rom[247] = 12'h000;
rom[248] = 12'h000;
rom[249] = 12'h000;
rom[250] = 12'h000;
rom[251] = 12'h000;
rom[252] = 12'h00f;
rom[253] = 12'h00f;
rom[254] = 12'h00f;
rom[255] = 12'h00f;
rom[256] = 12'h00f;
rom[257] = 12'h00f;
rom[258] = 12'h000;
rom[259] = 12'h000;
rom[260] = 12'h000;
rom[261] = 12'h000;
rom[262] = 12'h000;
rom[263] = 12'h000;
rom[264] = 12'h007;
rom[265] = 12'h007;
rom[266] = 12'h000;
rom[267] = 12'h000;
rom[268] = 12'h000;
rom[269] = 12'h000;
rom[270] = 12'h000;
rom[271] = 12'h000;
rom[272] = 12'h000;
rom[273] = 12'h000;
rom[274] = 12'h000;
rom[275] = 12'h000;
rom[276] = 12'h000;
rom[277] = 12'h000;
rom[278] = 12'h00f;
rom[279] = 12'h00f;
rom[280] = 12'h00f;
rom[281] = 12'h00f;
rom[282] = 12'h00f;
rom[283] = 12'h00f;
rom[284] = 12'h000;
rom[285] = 12'h000;
rom[286] = 12'h000;
rom[287] = 12'h000;
rom[288] = 12'h000;
rom[289] = 12'h000;
rom[290] = 12'h007;
rom[291] = 12'h007;
rom[292] = 12'h000;
rom[293] = 12'h000;
rom[294] = 12'h000;
rom[295] = 12'h000;
rom[296] = 12'h000;
rom[297] = 12'h000;
rom[298] = 12'h000;
rom[299] = 12'h000;
rom[300] = 12'h000;
rom[301] = 12'h000;
rom[302] = 12'h000;
rom[303] = 12'h000;
rom[304] = 12'h00f;
rom[305] = 12'h00f;
rom[306] = 12'h00f;
rom[307] = 12'h00f;
rom[308] = 12'h00f;
rom[309] = 12'h00f;
rom[310] = 12'h000;
rom[311] = 12'h000;
rom[312] = 12'h000;
rom[313] = 12'h000;
rom[314] = 12'h007;
rom[315] = 12'h007;
rom[316] = 12'h000;
rom[317] = 12'h000;
rom[318] = 12'h007;
rom[319] = 12'h007;
rom[320] = 12'h000;
rom[321] = 12'h000;
rom[322] = 12'h000;
rom[323] = 12'h000;
rom[324] = 12'h000;
rom[325] = 12'h000;
rom[326] = 12'h000;
rom[327] = 12'h000;
rom[328] = 12'h000;
rom[329] = 12'h000;
rom[330] = 12'h00f;
rom[331] = 12'h00f;
rom[332] = 12'h00f;
rom[333] = 12'h00f;
rom[334] = 12'h00f;
rom[335] = 12'h00f;
rom[336] = 12'h000;
rom[337] = 12'h000;
rom[338] = 12'h000;
rom[339] = 12'h000;
rom[340] = 12'h007;
rom[341] = 12'h007;
rom[342] = 12'h000;
rom[343] = 12'h000;
rom[344] = 12'h007;
rom[345] = 12'h007;
rom[346] = 12'h000;
rom[347] = 12'h000;
rom[348] = 12'h000;
rom[349] = 12'h000;
rom[350] = 12'h000;
rom[351] = 12'h000;
rom[352] = 12'h000;
rom[353] = 12'h000;
rom[354] = 12'h000;
rom[355] = 12'h000;
rom[356] = 12'h00f;
rom[357] = 12'h00f;
rom[358] = 12'h00f;
rom[359] = 12'h00f;
rom[360] = 12'h00f;
rom[361] = 12'h00f;
rom[362] = 12'h000;
rom[363] = 12'h000;
rom[364] = 12'h000;
rom[365] = 12'h000;
rom[366] = 12'h000;
rom[367] = 12'h000;
rom[368] = 12'h007;
rom[369] = 12'h007;
rom[370] = 12'h000;
rom[371] = 12'h000;
rom[372] = 12'h000;
rom[373] = 12'h000;
rom[374] = 12'h000;
rom[375] = 12'h000;
rom[376] = 12'h000;
rom[377] = 12'h000;
rom[378] = 12'h000;
rom[379] = 12'h000;
rom[380] = 12'h000;
rom[381] = 12'h000;
rom[382] = 12'h00f;
rom[383] = 12'h00f;
rom[384] = 12'h00f;
rom[385] = 12'h00f;
rom[386] = 12'h00f;
rom[387] = 12'h00f;
rom[388] = 12'h000;
rom[389] = 12'h000;
rom[390] = 12'h000;
rom[391] = 12'h000;
rom[392] = 12'h000;
rom[393] = 12'h000;
rom[394] = 12'h007;
rom[395] = 12'h007;
rom[396] = 12'h000;
rom[397] = 12'h000;
rom[398] = 12'h000;
rom[399] = 12'h000;
rom[400] = 12'h000;
rom[401] = 12'h000;
rom[402] = 12'h000;
rom[403] = 12'h000;
rom[404] = 12'h000;
rom[405] = 12'h000;
rom[406] = 12'h000;
rom[407] = 12'h000;
rom[408] = 12'h00f;
rom[409] = 12'h00f;
rom[410] = 12'h00f;
rom[411] = 12'h00f;
rom[412] = 12'h00f;
rom[413] = 12'h00f;
rom[414] = 12'h000;
rom[415] = 12'h000;
rom[416] = 12'h000;
rom[417] = 12'h000;
rom[418] = 12'h007;
rom[419] = 12'h007;
rom[420] = 12'h000;
rom[421] = 12'h000;
rom[422] = 12'h007;
rom[423] = 12'h007;
rom[424] = 12'h000;
rom[425] = 12'h000;
rom[426] = 12'h000;
rom[427] = 12'h000;
rom[428] = 12'h000;
rom[429] = 12'h000;
rom[430] = 12'h000;
rom[431] = 12'h000;
rom[432] = 12'h000;
rom[433] = 12'h000;
rom[434] = 12'h00f;
rom[435] = 12'h00f;
rom[436] = 12'h00f;
rom[437] = 12'h00f;
rom[438] = 12'h00f;
rom[439] = 12'h00f;
rom[440] = 12'h000;
rom[441] = 12'h000;
rom[442] = 12'h000;
rom[443] = 12'h000;
rom[444] = 12'h007;
rom[445] = 12'h007;
rom[446] = 12'h000;
rom[447] = 12'h000;
rom[448] = 12'h007;
rom[449] = 12'h007;
rom[450] = 12'h000;
rom[451] = 12'h000;
rom[452] = 12'h000;
rom[453] = 12'h000;
rom[454] = 12'h000;
rom[455] = 12'h000;
rom[456] = 12'h000;
rom[457] = 12'h000;
rom[458] = 12'h000;
rom[459] = 12'h000;
rom[460] = 12'h00f;
rom[461] = 12'h00f;
rom[462] = 12'h00f;
rom[463] = 12'h00f;
rom[464] = 12'h00f;
rom[465] = 12'h00f;
rom[466] = 12'h000;
rom[467] = 12'h000;
rom[468] = 12'h000;
rom[469] = 12'h000;
rom[470] = 12'h000;
rom[471] = 12'h000;
rom[472] = 12'h007;
rom[473] = 12'h007;
rom[474] = 12'h000;
rom[475] = 12'h000;
rom[476] = 12'h000;
rom[477] = 12'h000;
rom[478] = 12'h000;
rom[479] = 12'h000;
rom[480] = 12'h000;
rom[481] = 12'h000;
rom[482] = 12'h000;
rom[483] = 12'h000;
rom[484] = 12'h000;
rom[485] = 12'h000;
rom[486] = 12'h000;
rom[487] = 12'h000;
rom[488] = 12'h00f;
rom[489] = 12'h00f;
rom[490] = 12'h00f;
rom[491] = 12'h00f;
rom[492] = 12'h000;
rom[493] = 12'h000;
rom[494] = 12'h000;
rom[495] = 12'h000;
rom[496] = 12'h000;
rom[497] = 12'h000;
rom[498] = 12'h007;
rom[499] = 12'h007;
rom[500] = 12'h000;
rom[501] = 12'h000;
rom[502] = 12'h000;
rom[503] = 12'h000;
rom[504] = 12'h000;
rom[505] = 12'h000;
rom[506] = 12'h000;
rom[507] = 12'h000;
rom[508] = 12'h000;
rom[509] = 12'h000;
rom[510] = 12'h000;
rom[511] = 12'h000;
rom[512] = 12'h000;
rom[513] = 12'h000;
rom[514] = 12'h00f;
rom[515] = 12'h00f;
rom[516] = 12'h00f;
rom[517] = 12'h00f;
rom[518] = 12'h000;
rom[519] = 12'h000;
rom[520] = 12'h000;
rom[521] = 12'h000;
rom[522] = 12'h007;
rom[523] = 12'h007;
rom[524] = 12'h000;
rom[525] = 12'h000;
rom[526] = 12'h000;
rom[527] = 12'h000;
rom[528] = 12'h007;
rom[529] = 12'h007;
rom[530] = 12'h000;
rom[531] = 12'h000;
rom[532] = 12'h007;
rom[533] = 12'h007;
rom[534] = 12'h000;
rom[535] = 12'h000;
rom[536] = 12'h007;
rom[537] = 12'h007;
rom[538] = 12'h000;
rom[539] = 12'h000;
rom[540] = 12'h000;
rom[541] = 12'h000;
rom[542] = 12'h00f;
rom[543] = 12'h00f;
rom[544] = 12'h000;
rom[545] = 12'h000;
rom[546] = 12'h000;
rom[547] = 12'h000;
rom[548] = 12'h007;
rom[549] = 12'h007;
rom[550] = 12'h000;
rom[551] = 12'h000;
rom[552] = 12'h000;
rom[553] = 12'h000;
rom[554] = 12'h007;
rom[555] = 12'h007;
rom[556] = 12'h000;
rom[557] = 12'h000;
rom[558] = 12'h007;
rom[559] = 12'h007;
rom[560] = 12'h000;
rom[561] = 12'h000;
rom[562] = 12'h007;
rom[563] = 12'h007;
rom[564] = 12'h000;
rom[565] = 12'h000;
rom[566] = 12'h000;
rom[567] = 12'h000;
rom[568] = 12'h00f;
rom[569] = 12'h00f;
rom[570] = 12'h000;
rom[571] = 12'h000;
rom[572] = 12'h000;
rom[573] = 12'h000;
rom[574] = 12'h000;
rom[575] = 12'h000;
rom[576] = 12'h000;
rom[577] = 12'h000;
rom[578] = 12'h007;
rom[579] = 12'h007;
rom[580] = 12'h000;
rom[581] = 12'h000;
rom[582] = 12'h007;
rom[583] = 12'h007;
rom[584] = 12'h000;
rom[585] = 12'h000;
rom[586] = 12'h007;
rom[587] = 12'h007;
rom[588] = 12'h000;
rom[589] = 12'h000;
rom[590] = 12'h007;
rom[591] = 12'h007;
rom[592] = 12'h000;
rom[593] = 12'h000;
rom[594] = 12'h000;
rom[595] = 12'h000;
rom[596] = 12'h000;
rom[597] = 12'h000;
rom[598] = 12'h000;
rom[599] = 12'h000;
rom[600] = 12'h000;
rom[601] = 12'h000;
rom[602] = 12'h000;
rom[603] = 12'h000;
rom[604] = 12'h007;
rom[605] = 12'h007;
rom[606] = 12'h000;
rom[607] = 12'h000;
rom[608] = 12'h007;
rom[609] = 12'h007;
rom[610] = 12'h000;
rom[611] = 12'h000;
rom[612] = 12'h007;
rom[613] = 12'h007;
rom[614] = 12'h000;
rom[615] = 12'h000;
rom[616] = 12'h007;
rom[617] = 12'h007;
rom[618] = 12'h000;
rom[619] = 12'h000;
rom[620] = 12'h000;
rom[621] = 12'h000;
rom[622] = 12'h000;
rom[623] = 12'h000;
rom[624] = 12'h000;
rom[625] = 12'h000;
rom[626] = 12'h007;
rom[627] = 12'h007;
rom[628] = 12'h000;
rom[629] = 12'h000;
rom[630] = 12'h000;
rom[631] = 12'h000;
rom[632] = 12'h007;
rom[633] = 12'h007;
rom[634] = 12'h000;
rom[635] = 12'h000;
rom[636] = 12'h007;
rom[637] = 12'h007;
rom[638] = 12'h000;
rom[639] = 12'h000;
rom[640] = 12'h007;
rom[641] = 12'h007;
rom[642] = 12'h000;
rom[643] = 12'h000;
rom[644] = 12'h000;
rom[645] = 12'h000;
rom[646] = 12'h00f;
rom[647] = 12'h00f;
rom[648] = 12'h000;
rom[649] = 12'h000;
rom[650] = 12'h000;
rom[651] = 12'h000;
rom[652] = 12'h007;
rom[653] = 12'h007;
rom[654] = 12'h000;
rom[655] = 12'h000;
rom[656] = 12'h000;
rom[657] = 12'h000;
rom[658] = 12'h007;
rom[659] = 12'h007;
rom[660] = 12'h000;
rom[661] = 12'h000;
rom[662] = 12'h007;
rom[663] = 12'h007;
rom[664] = 12'h000;
rom[665] = 12'h000;
rom[666] = 12'h007;
rom[667] = 12'h007;
rom[668] = 12'h000;
rom[669] = 12'h000;
rom[670] = 12'h000;
rom[671] = 12'h000;
rom[672] = 12'h00f;
rom[673] = 12'h00f;
rom[674] = 12'h000;
rom[675] = 12'h000;
rom[676] = 12'h000;
rom[677] = 12'h000;
rom[678] = 12'h000;
rom[679] = 12'h000;
rom[680] = 12'h007;
rom[681] = 12'h007;
rom[682] = 12'h000;
rom[683] = 12'h000;
rom[684] = 12'h000;
rom[685] = 12'h000;
rom[686] = 12'h000;
rom[687] = 12'h000;
rom[688] = 12'h000;
rom[689] = 12'h000;
rom[690] = 12'h000;
rom[691] = 12'h000;
rom[692] = 12'h000;
rom[693] = 12'h000;
rom[694] = 12'h000;
rom[695] = 12'h000;
rom[696] = 12'h00f;
rom[697] = 12'h00f;
rom[698] = 12'h00f;
rom[699] = 12'h00f;
rom[700] = 12'h000;
rom[701] = 12'h000;
rom[702] = 12'h000;
rom[703] = 12'h000;
rom[704] = 12'h000;
rom[705] = 12'h000;
rom[706] = 12'h007;
rom[707] = 12'h007;
rom[708] = 12'h000;
rom[709] = 12'h000;
rom[710] = 12'h000;
rom[711] = 12'h000;
rom[712] = 12'h000;
rom[713] = 12'h000;
rom[714] = 12'h000;
rom[715] = 12'h000;
rom[716] = 12'h000;
rom[717] = 12'h000;
rom[718] = 12'h000;
rom[719] = 12'h000;
rom[720] = 12'h000;
rom[721] = 12'h000;
rom[722] = 12'h00f;
rom[723] = 12'h00f;
rom[724] = 12'h00f;
rom[725] = 12'h00f;
rom[726] = 12'h000;
rom[727] = 12'h000;
rom[728] = 12'h000;
rom[729] = 12'h000;
rom[730] = 12'h007;
rom[731] = 12'h007;
rom[732] = 12'h000;
rom[733] = 12'h000;
rom[734] = 12'h007;
rom[735] = 12'h007;
rom[736] = 12'h000;
rom[737] = 12'h000;
rom[738] = 12'h000;
rom[739] = 12'h000;
rom[740] = 12'h000;
rom[741] = 12'h000;
rom[742] = 12'h000;
rom[743] = 12'h000;
rom[744] = 12'h000;
rom[745] = 12'h000;
rom[746] = 12'h00f;
rom[747] = 12'h00f;
rom[748] = 12'h00f;
rom[749] = 12'h00f;
rom[750] = 12'h00f;
rom[751] = 12'h00f;
rom[752] = 12'h000;
rom[753] = 12'h000;
rom[754] = 12'h000;
rom[755] = 12'h000;
rom[756] = 12'h007;
rom[757] = 12'h007;
rom[758] = 12'h000;
rom[759] = 12'h000;
rom[760] = 12'h007;
rom[761] = 12'h007;
rom[762] = 12'h000;
rom[763] = 12'h000;
rom[764] = 12'h000;
rom[765] = 12'h000;
rom[766] = 12'h000;
rom[767] = 12'h000;
rom[768] = 12'h000;
rom[769] = 12'h000;
rom[770] = 12'h000;
rom[771] = 12'h000;
rom[772] = 12'h00f;
rom[773] = 12'h00f;
rom[774] = 12'h00f;
rom[775] = 12'h00f;
rom[776] = 12'h00f;
rom[777] = 12'h00f;
rom[778] = 12'h000;
rom[779] = 12'h000;
rom[780] = 12'h000;
rom[781] = 12'h000;
rom[782] = 12'h000;
rom[783] = 12'h000;
rom[784] = 12'h007;
rom[785] = 12'h007;
rom[786] = 12'h000;
rom[787] = 12'h000;
rom[788] = 12'h000;
rom[789] = 12'h000;
rom[790] = 12'h000;
rom[791] = 12'h000;
rom[792] = 12'h000;
rom[793] = 12'h000;
rom[794] = 12'h000;
rom[795] = 12'h000;
rom[796] = 12'h000;
rom[797] = 12'h000;
rom[798] = 12'h00f;
rom[799] = 12'h00f;
rom[800] = 12'h00f;
rom[801] = 12'h00f;
rom[802] = 12'h00f;
rom[803] = 12'h00f;
rom[804] = 12'h000;
rom[805] = 12'h000;
rom[806] = 12'h000;
rom[807] = 12'h000;
rom[808] = 12'h000;
rom[809] = 12'h000;
rom[810] = 12'h007;
rom[811] = 12'h007;
rom[812] = 12'h000;
rom[813] = 12'h000;
rom[814] = 12'h000;
rom[815] = 12'h000;
rom[816] = 12'h000;
rom[817] = 12'h000;
rom[818] = 12'h000;
rom[819] = 12'h000;
rom[820] = 12'h000;
rom[821] = 12'h000;
rom[822] = 12'h000;
rom[823] = 12'h000;
rom[824] = 12'h00f;
rom[825] = 12'h00f;
rom[826] = 12'h00f;
rom[827] = 12'h00f;
rom[828] = 12'h00f;
rom[829] = 12'h00f;
rom[830] = 12'h000;
rom[831] = 12'h000;
rom[832] = 12'h000;
rom[833] = 12'h000;
rom[834] = 12'h007;
rom[835] = 12'h007;
rom[836] = 12'h000;
rom[837] = 12'h000;
rom[838] = 12'h007;
rom[839] = 12'h007;
rom[840] = 12'h000;
rom[841] = 12'h000;
rom[842] = 12'h000;
rom[843] = 12'h000;
rom[844] = 12'h000;
rom[845] = 12'h000;
rom[846] = 12'h000;
rom[847] = 12'h000;
rom[848] = 12'h000;
rom[849] = 12'h000;
rom[850] = 12'h00f;
rom[851] = 12'h00f;
rom[852] = 12'h00f;
rom[853] = 12'h00f;
rom[854] = 12'h00f;
rom[855] = 12'h00f;
rom[856] = 12'h000;
rom[857] = 12'h000;
rom[858] = 12'h000;
rom[859] = 12'h000;
rom[860] = 12'h007;
rom[861] = 12'h007;
rom[862] = 12'h000;
rom[863] = 12'h000;
rom[864] = 12'h007;
rom[865] = 12'h007;
rom[866] = 12'h000;
rom[867] = 12'h000;
rom[868] = 12'h000;
rom[869] = 12'h000;
rom[870] = 12'h000;
rom[871] = 12'h000;
rom[872] = 12'h000;
rom[873] = 12'h000;
rom[874] = 12'h000;
rom[875] = 12'h000;
rom[876] = 12'h00f;
rom[877] = 12'h00f;
rom[878] = 12'h00f;
rom[879] = 12'h00f;
rom[880] = 12'h00f;
rom[881] = 12'h00f;
rom[882] = 12'h000;
rom[883] = 12'h000;
rom[884] = 12'h000;
rom[885] = 12'h000;
rom[886] = 12'h000;
rom[887] = 12'h000;
rom[888] = 12'h007;
rom[889] = 12'h007;
rom[890] = 12'h000;
rom[891] = 12'h000;
rom[892] = 12'h000;
rom[893] = 12'h000;
rom[894] = 12'h000;
rom[895] = 12'h000;
rom[896] = 12'h000;
rom[897] = 12'h000;
rom[898] = 12'h000;
rom[899] = 12'h000;
rom[900] = 12'h000;
rom[901] = 12'h000;
rom[902] = 12'h00f;
rom[903] = 12'h00f;
rom[904] = 12'h00f;
rom[905] = 12'h00f;
rom[906] = 12'h00f;
rom[907] = 12'h00f;
rom[908] = 12'h000;
rom[909] = 12'h000;
rom[910] = 12'h000;
rom[911] = 12'h000;
rom[912] = 12'h000;
rom[913] = 12'h000;
rom[914] = 12'h007;
rom[915] = 12'h007;
rom[916] = 12'h000;
rom[917] = 12'h000;
rom[918] = 12'h000;
rom[919] = 12'h000;
rom[920] = 12'h000;
rom[921] = 12'h000;
rom[922] = 12'h000;
rom[923] = 12'h000;
rom[924] = 12'h000;
rom[925] = 12'h000;
rom[926] = 12'h000;
rom[927] = 12'h000;
rom[928] = 12'h00f;
rom[929] = 12'h00f;
rom[930] = 12'h00f;
rom[931] = 12'h00f;
rom[932] = 12'h00f;
rom[933] = 12'h00f;
rom[934] = 12'h000;
rom[935] = 12'h000;
rom[936] = 12'h000;
rom[937] = 12'h000;
rom[938] = 12'h007;
rom[939] = 12'h007;
rom[940] = 12'h000;
rom[941] = 12'h000;
rom[942] = 12'h007;
rom[943] = 12'h007;
rom[944] = 12'h000;
rom[945] = 12'h000;
rom[946] = 12'h000;
rom[947] = 12'h000;
rom[948] = 12'h000;
rom[949] = 12'h000;
rom[950] = 12'h000;
rom[951] = 12'h000;
rom[952] = 12'h000;
rom[953] = 12'h000;
rom[954] = 12'h00f;
rom[955] = 12'h00f;
rom[956] = 12'h00f;
rom[957] = 12'h00f;
rom[958] = 12'h00f;
rom[959] = 12'h00f;
rom[960] = 12'h000;
rom[961] = 12'h000;
rom[962] = 12'h000;
rom[963] = 12'h000;
rom[964] = 12'h007;
rom[965] = 12'h007;
rom[966] = 12'h000;
rom[967] = 12'h000;
rom[968] = 12'h007;
rom[969] = 12'h007;
rom[970] = 12'h000;
rom[971] = 12'h000;
rom[972] = 12'h000;
rom[973] = 12'h000;
rom[974] = 12'h000;
rom[975] = 12'h000;
rom[976] = 12'h000;
rom[977] = 12'h000;
rom[978] = 12'h000;
rom[979] = 12'h000;
rom[980] = 12'h00f;
rom[981] = 12'h00f;
rom[982] = 12'h00f;
rom[983] = 12'h00f;
rom[984] = 12'h00f;
rom[985] = 12'h00f;
rom[986] = 12'h000;
rom[987] = 12'h000;
rom[988] = 12'h000;
rom[989] = 12'h000;
rom[990] = 12'h000;
rom[991] = 12'h000;
rom[992] = 12'h007;
rom[993] = 12'h007;
rom[994] = 12'h000;
rom[995] = 12'h000;
rom[996] = 12'h000;
rom[997] = 12'h000;
rom[998] = 12'h007;
rom[999] = 12'h007;
rom[1000] = 12'h000;
rom[1001] = 12'h000;
rom[1002] = 12'h007;
rom[1003] = 12'h007;
rom[1004] = 12'h000;
rom[1005] = 12'h000;
rom[1006] = 12'h000;
rom[1007] = 12'h000;
rom[1008] = 12'h00f;
rom[1009] = 12'h00f;
rom[1010] = 12'h00f;
rom[1011] = 12'h00f;
rom[1012] = 12'h000;
rom[1013] = 12'h000;
rom[1014] = 12'h000;
rom[1015] = 12'h000;
rom[1016] = 12'h000;
rom[1017] = 12'h000;
rom[1018] = 12'h007;
rom[1019] = 12'h007;
rom[1020] = 12'h000;
rom[1021] = 12'h000;
rom[1022] = 12'h000;
rom[1023] = 12'h000;
rom[1024] = 12'h007;
rom[1025] = 12'h007;
rom[1026] = 12'h000;
rom[1027] = 12'h000;
rom[1028] = 12'h007;
rom[1029] = 12'h007;
rom[1030] = 12'h000;
rom[1031] = 12'h000;
rom[1032] = 12'h000;
rom[1033] = 12'h000;
rom[1034] = 12'h00f;
rom[1035] = 12'h00f;
rom[1036] = 12'h00f;
rom[1037] = 12'h00f;
rom[1038] = 12'h000;
rom[1039] = 12'h000;
rom[1040] = 12'h000;
rom[1041] = 12'h000;
rom[1042] = 12'h007;
rom[1043] = 12'h007;
rom[1044] = 12'h000;
rom[1045] = 12'h000;
rom[1046] = 12'h000;
rom[1047] = 12'h000;
rom[1048] = 12'h007;
rom[1049] = 12'h007;
rom[1050] = 12'h000;
rom[1051] = 12'h000;
rom[1052] = 12'h007;
rom[1053] = 12'h007;
rom[1054] = 12'h000;
rom[1055] = 12'h000;
rom[1056] = 12'h007;
rom[1057] = 12'h007;
rom[1058] = 12'h000;
rom[1059] = 12'h000;
rom[1060] = 12'h000;
rom[1061] = 12'h000;
rom[1062] = 12'h00f;
rom[1063] = 12'h00f;
rom[1064] = 12'h000;
rom[1065] = 12'h000;
rom[1066] = 12'h000;
rom[1067] = 12'h000;
rom[1068] = 12'h007;
rom[1069] = 12'h007;
rom[1070] = 12'h000;
rom[1071] = 12'h000;
rom[1072] = 12'h000;
rom[1073] = 12'h000;
rom[1074] = 12'h007;
rom[1075] = 12'h007;
rom[1076] = 12'h000;
rom[1077] = 12'h000;
rom[1078] = 12'h007;
rom[1079] = 12'h007;
rom[1080] = 12'h000;
rom[1081] = 12'h000;
rom[1082] = 12'h007;
rom[1083] = 12'h007;
rom[1084] = 12'h000;
rom[1085] = 12'h000;
rom[1086] = 12'h000;
rom[1087] = 12'h000;
rom[1088] = 12'h00f;
rom[1089] = 12'h00f;
rom[1090] = 12'h000;
rom[1091] = 12'h000;
rom[1092] = 12'h000;
rom[1093] = 12'h000;
rom[1094] = 12'h000;
rom[1095] = 12'h000;
rom[1096] = 12'h000;
rom[1097] = 12'h000;
rom[1098] = 12'h007;
rom[1099] = 12'h007;
rom[1100] = 12'h000;
rom[1101] = 12'h000;
rom[1102] = 12'h007;
rom[1103] = 12'h007;
rom[1104] = 12'h000;
rom[1105] = 12'h000;
rom[1106] = 12'h007;
rom[1107] = 12'h007;
rom[1108] = 12'h000;
rom[1109] = 12'h000;
rom[1110] = 12'h007;
rom[1111] = 12'h007;
rom[1112] = 12'h000;
rom[1113] = 12'h000;
rom[1114] = 12'h000;
rom[1115] = 12'h000;
rom[1116] = 12'h000;
rom[1117] = 12'h000;
rom[1118] = 12'h000;
rom[1119] = 12'h000;
rom[1120] = 12'h000;
rom[1121] = 12'h000;
rom[1122] = 12'h000;
rom[1123] = 12'h000;
rom[1124] = 12'h007;
rom[1125] = 12'h007;
rom[1126] = 12'h000;
rom[1127] = 12'h000;
rom[1128] = 12'h007;
rom[1129] = 12'h007;
rom[1130] = 12'h000;
rom[1131] = 12'h000;
rom[1132] = 12'h007;
rom[1133] = 12'h007;
rom[1134] = 12'h000;
rom[1135] = 12'h000;
rom[1136] = 12'h007;
rom[1137] = 12'h007;
rom[1138] = 12'h000;
rom[1139] = 12'h000;
rom[1140] = 12'h000;
rom[1141] = 12'h000;
rom[1142] = 12'h000;
rom[1143] = 12'h000;
rom[1144] = 12'h000;
rom[1145] = 12'h000;
rom[1146] = 12'h000;
rom[1147] = 12'h000;
rom[1148] = 12'h000;
rom[1149] = 12'h000;
rom[1150] = 12'h000;
rom[1151] = 12'h000;
rom[1152] = 12'h000;
rom[1153] = 12'h000;
rom[1154] = 12'h000;
rom[1155] = 12'h000;
rom[1156] = 12'h000;
rom[1157] = 12'h000;
rom[1158] = 12'h000;
rom[1159] = 12'h000;
rom[1160] = 12'h000;
rom[1161] = 12'h000;
rom[1162] = 12'h000;
rom[1163] = 12'h000;
rom[1164] = 12'h000;
rom[1165] = 12'h000;
rom[1166] = 12'h000;
rom[1167] = 12'h000;
rom[1168] = 12'h000;
rom[1169] = 12'h000;
rom[1170] = 12'h000;
rom[1171] = 12'h000;
rom[1172] = 12'h000;
rom[1173] = 12'h000;
rom[1174] = 12'h000;
rom[1175] = 12'h000;
rom[1176] = 12'h000;
rom[1177] = 12'h000;
rom[1178] = 12'h000;
rom[1179] = 12'h000;
rom[1180] = 12'h000;
rom[1181] = 12'h000;
rom[1182] = 12'h000;
rom[1183] = 12'h000;
rom[1184] = 12'h000;
rom[1185] = 12'h000;
rom[1186] = 12'h000;
rom[1187] = 12'h000;
rom[1188] = 12'h000;
rom[1189] = 12'h000;
rom[1190] = 12'h000;
rom[1191] = 12'h000;
rom[1192] = 12'h000;
rom[1193] = 12'h000;
rom[1194] = 12'h000;
rom[1195] = 12'h000;

  end
  endmodule

    module dash_rom (                       //восемь
  input  wire    [13:0]     addr,
  output wire    [11:0]     word
);

  logic [11:0] rom [(46 * 26)];

  assign word = rom[addr];

  initial begin
rom[0] = 12'h000;
rom[1] = 12'h000;
rom[2] = 12'h000;
rom[3] = 12'h000;
rom[4] = 12'h000;
rom[5] = 12'h000;
rom[6] = 12'h000;
rom[7] = 12'h000;
rom[8] = 12'h000;
rom[9] = 12'h000;
rom[10] = 12'h000;
rom[11] = 12'h000;
rom[12] = 12'h000;
rom[13] = 12'h000;
rom[14] = 12'h000;
rom[15] = 12'h000;
rom[16] = 12'h000;
rom[17] = 12'h000;
rom[18] = 12'h000;
rom[19] = 12'h000;
rom[20] = 12'h000;
rom[21] = 12'h000;
rom[22] = 12'h000;
rom[23] = 12'h000;
rom[24] = 12'h000;
rom[25] = 12'h000;
rom[26] = 12'h000;
rom[27] = 12'h000;
rom[28] = 12'h000;
rom[29] = 12'h000;
rom[30] = 12'h000;
rom[31] = 12'h000;
rom[32] = 12'h000;
rom[33] = 12'h000;
rom[34] = 12'h000;
rom[35] = 12'h000;
rom[36] = 12'h000;
rom[37] = 12'h000;
rom[38] = 12'h000;
rom[39] = 12'h000;
rom[40] = 12'h000;
rom[41] = 12'h000;
rom[42] = 12'h000;
rom[43] = 12'h000;
rom[44] = 12'h000;
rom[45] = 12'h000;
rom[46] = 12'h000;
rom[47] = 12'h000;
rom[48] = 12'h000;
rom[49] = 12'h000;
rom[50] = 12'h000;
rom[51] = 12'h000;
rom[52] = 12'h000;
rom[53] = 12'h000;
rom[54] = 12'h000;
rom[55] = 12'h000;
rom[56] = 12'h00f;
rom[57] = 12'h00f;
rom[58] = 12'h00f;
rom[59] = 12'h00f;
rom[60] = 12'h00f;
rom[61] = 12'h00f;
rom[62] = 12'h00f;
rom[63] = 12'h00f;
rom[64] = 12'h00f;
rom[65] = 12'h00f;
rom[66] = 12'h00f;
rom[67] = 12'h00f;
rom[68] = 12'h00f;
rom[69] = 12'h00f;
rom[70] = 12'h00f;
rom[71] = 12'h00f;
rom[72] = 12'h00f;
rom[73] = 12'h00f;
rom[74] = 12'h000;
rom[75] = 12'h000;
rom[76] = 12'h000;
rom[77] = 12'h000;
rom[78] = 12'h000;
rom[79] = 12'h000;
rom[80] = 12'h000;
rom[81] = 12'h000;
rom[82] = 12'h00f;
rom[83] = 12'h00f;
rom[84] = 12'h00f;
rom[85] = 12'h00f;
rom[86] = 12'h00f;
rom[87] = 12'h00f;
rom[88] = 12'h00f;
rom[89] = 12'h00f;
rom[90] = 12'h00f;
rom[91] = 12'h00f;
rom[92] = 12'h00f;
rom[93] = 12'h00f;
rom[94] = 12'h00f;
rom[95] = 12'h00f;
rom[96] = 12'h00f;
rom[97] = 12'h00f;
rom[98] = 12'h00f;
rom[99] = 12'h00f;
rom[100] = 12'h000;
rom[101] = 12'h000;
rom[102] = 12'h000;
rom[103] = 12'h000;
rom[104] = 12'h000;
rom[105] = 12'h000;
rom[106] = 12'h00f;
rom[107] = 12'h00f;
rom[108] = 12'h000;
rom[109] = 12'h000;
rom[110] = 12'h00f;
rom[111] = 12'h00f;
rom[112] = 12'h00f;
rom[113] = 12'h00f;
rom[114] = 12'h00f;
rom[115] = 12'h00f;
rom[116] = 12'h00f;
rom[117] = 12'h00f;
rom[118] = 12'h00f;
rom[119] = 12'h00f;
rom[120] = 12'h00f;
rom[121] = 12'h00f;
rom[122] = 12'h00f;
rom[123] = 12'h00f;
rom[124] = 12'h000;
rom[125] = 12'h000;
rom[126] = 12'h00f;
rom[127] = 12'h00f;
rom[128] = 12'h000;
rom[129] = 12'h000;
rom[130] = 12'h000;
rom[131] = 12'h000;
rom[132] = 12'h00f;
rom[133] = 12'h00f;
rom[134] = 12'h000;
rom[135] = 12'h000;
rom[136] = 12'h00f;
rom[137] = 12'h00f;
rom[138] = 12'h00f;
rom[139] = 12'h00f;
rom[140] = 12'h00f;
rom[141] = 12'h00f;
rom[142] = 12'h00f;
rom[143] = 12'h00f;
rom[144] = 12'h00f;
rom[145] = 12'h00f;
rom[146] = 12'h00f;
rom[147] = 12'h00f;
rom[148] = 12'h00f;
rom[149] = 12'h00f;
rom[150] = 12'h000;
rom[151] = 12'h000;
rom[152] = 12'h00f;
rom[153] = 12'h00f;
rom[154] = 12'h000;
rom[155] = 12'h000;
rom[156] = 12'h000;
rom[157] = 12'h000;
rom[158] = 12'h00f;
rom[159] = 12'h00f;
rom[160] = 12'h00f;
rom[161] = 12'h00f;
rom[162] = 12'h000;
rom[163] = 12'h000;
rom[164] = 12'h00f;
rom[165] = 12'h00f;
rom[166] = 12'h00f;
rom[167] = 12'h00f;
rom[168] = 12'h00f;
rom[169] = 12'h00f;
rom[170] = 12'h00f;
rom[171] = 12'h00f;
rom[172] = 12'h00f;
rom[173] = 12'h00f;
rom[174] = 12'h000;
rom[175] = 12'h000;
rom[176] = 12'h00f;
rom[177] = 12'h00f;
rom[178] = 12'h00f;
rom[179] = 12'h00f;
rom[180] = 12'h000;
rom[181] = 12'h000;
rom[182] = 12'h000;
rom[183] = 12'h000;
rom[184] = 12'h00f;
rom[185] = 12'h00f;
rom[186] = 12'h00f;
rom[187] = 12'h00f;
rom[188] = 12'h000;
rom[189] = 12'h000;
rom[190] = 12'h00f;
rom[191] = 12'h00f;
rom[192] = 12'h00f;
rom[193] = 12'h00f;
rom[194] = 12'h00f;
rom[195] = 12'h00f;
rom[196] = 12'h00f;
rom[197] = 12'h00f;
rom[198] = 12'h00f;
rom[199] = 12'h00f;
rom[200] = 12'h000;
rom[201] = 12'h000;
rom[202] = 12'h00f;
rom[203] = 12'h00f;
rom[204] = 12'h00f;
rom[205] = 12'h00f;
rom[206] = 12'h000;
rom[207] = 12'h000;
rom[208] = 12'h000;
rom[209] = 12'h000;
rom[210] = 12'h00f;
rom[211] = 12'h00f;
rom[212] = 12'h00f;
rom[213] = 12'h00f;
rom[214] = 12'h00f;
rom[215] = 12'h00f;
rom[216] = 12'h000;
rom[217] = 12'h000;
rom[218] = 12'h000;
rom[219] = 12'h000;
rom[220] = 12'h000;
rom[221] = 12'h000;
rom[222] = 12'h000;
rom[223] = 12'h000;
rom[224] = 12'h000;
rom[225] = 12'h000;
rom[226] = 12'h00f;
rom[227] = 12'h00f;
rom[228] = 12'h00f;
rom[229] = 12'h00f;
rom[230] = 12'h00f;
rom[231] = 12'h00f;
rom[232] = 12'h000;
rom[233] = 12'h000;
rom[234] = 12'h000;
rom[235] = 12'h000;
rom[236] = 12'h00f;
rom[237] = 12'h00f;
rom[238] = 12'h00f;
rom[239] = 12'h00f;
rom[240] = 12'h00f;
rom[241] = 12'h00f;
rom[242] = 12'h000;
rom[243] = 12'h000;
rom[244] = 12'h000;
rom[245] = 12'h000;
rom[246] = 12'h000;
rom[247] = 12'h000;
rom[248] = 12'h000;
rom[249] = 12'h000;
rom[250] = 12'h000;
rom[251] = 12'h000;
rom[252] = 12'h00f;
rom[253] = 12'h00f;
rom[254] = 12'h00f;
rom[255] = 12'h00f;
rom[256] = 12'h00f;
rom[257] = 12'h00f;
rom[258] = 12'h000;
rom[259] = 12'h000;
rom[260] = 12'h000;
rom[261] = 12'h000;
rom[262] = 12'h00f;
rom[263] = 12'h00f;
rom[264] = 12'h00f;
rom[265] = 12'h00f;
rom[266] = 12'h00f;
rom[267] = 12'h00f;
rom[268] = 12'h000;
rom[269] = 12'h000;
rom[270] = 12'h000;
rom[271] = 12'h000;
rom[272] = 12'h000;
rom[273] = 12'h000;
rom[274] = 12'h000;
rom[275] = 12'h000;
rom[276] = 12'h000;
rom[277] = 12'h000;
rom[278] = 12'h00f;
rom[279] = 12'h00f;
rom[280] = 12'h00f;
rom[281] = 12'h00f;
rom[282] = 12'h00f;
rom[283] = 12'h00f;
rom[284] = 12'h000;
rom[285] = 12'h000;
rom[286] = 12'h000;
rom[287] = 12'h000;
rom[288] = 12'h00f;
rom[289] = 12'h00f;
rom[290] = 12'h00f;
rom[291] = 12'h00f;
rom[292] = 12'h00f;
rom[293] = 12'h00f;
rom[294] = 12'h000;
rom[295] = 12'h000;
rom[296] = 12'h000;
rom[297] = 12'h000;
rom[298] = 12'h000;
rom[299] = 12'h000;
rom[300] = 12'h000;
rom[301] = 12'h000;
rom[302] = 12'h000;
rom[303] = 12'h000;
rom[304] = 12'h00f;
rom[305] = 12'h00f;
rom[306] = 12'h00f;
rom[307] = 12'h00f;
rom[308] = 12'h00f;
rom[309] = 12'h00f;
rom[310] = 12'h000;
rom[311] = 12'h000;
rom[312] = 12'h000;
rom[313] = 12'h000;
rom[314] = 12'h00f;
rom[315] = 12'h00f;
rom[316] = 12'h00f;
rom[317] = 12'h00f;
rom[318] = 12'h00f;
rom[319] = 12'h00f;
rom[320] = 12'h000;
rom[321] = 12'h000;
rom[322] = 12'h000;
rom[323] = 12'h000;
rom[324] = 12'h000;
rom[325] = 12'h000;
rom[326] = 12'h000;
rom[327] = 12'h000;
rom[328] = 12'h000;
rom[329] = 12'h000;
rom[330] = 12'h00f;
rom[331] = 12'h00f;
rom[332] = 12'h00f;
rom[333] = 12'h00f;
rom[334] = 12'h00f;
rom[335] = 12'h00f;
rom[336] = 12'h000;
rom[337] = 12'h000;
rom[338] = 12'h000;
rom[339] = 12'h000;
rom[340] = 12'h00f;
rom[341] = 12'h00f;
rom[342] = 12'h00f;
rom[343] = 12'h00f;
rom[344] = 12'h00f;
rom[345] = 12'h00f;
rom[346] = 12'h000;
rom[347] = 12'h000;
rom[348] = 12'h000;
rom[349] = 12'h000;
rom[350] = 12'h000;
rom[351] = 12'h000;
rom[352] = 12'h000;
rom[353] = 12'h000;
rom[354] = 12'h000;
rom[355] = 12'h000;
rom[356] = 12'h00f;
rom[357] = 12'h00f;
rom[358] = 12'h00f;
rom[359] = 12'h00f;
rom[360] = 12'h00f;
rom[361] = 12'h00f;
rom[362] = 12'h000;
rom[363] = 12'h000;
rom[364] = 12'h000;
rom[365] = 12'h000;
rom[366] = 12'h00f;
rom[367] = 12'h00f;
rom[368] = 12'h00f;
rom[369] = 12'h00f;
rom[370] = 12'h00f;
rom[371] = 12'h00f;
rom[372] = 12'h000;
rom[373] = 12'h000;
rom[374] = 12'h000;
rom[375] = 12'h000;
rom[376] = 12'h000;
rom[377] = 12'h000;
rom[378] = 12'h000;
rom[379] = 12'h000;
rom[380] = 12'h000;
rom[381] = 12'h000;
rom[382] = 12'h00f;
rom[383] = 12'h00f;
rom[384] = 12'h00f;
rom[385] = 12'h00f;
rom[386] = 12'h00f;
rom[387] = 12'h00f;
rom[388] = 12'h000;
rom[389] = 12'h000;
rom[390] = 12'h000;
rom[391] = 12'h000;
rom[392] = 12'h00f;
rom[393] = 12'h00f;
rom[394] = 12'h00f;
rom[395] = 12'h00f;
rom[396] = 12'h00f;
rom[397] = 12'h00f;
rom[398] = 12'h000;
rom[399] = 12'h000;
rom[400] = 12'h000;
rom[401] = 12'h000;
rom[402] = 12'h000;
rom[403] = 12'h000;
rom[404] = 12'h000;
rom[405] = 12'h000;
rom[406] = 12'h000;
rom[407] = 12'h000;
rom[408] = 12'h00f;
rom[409] = 12'h00f;
rom[410] = 12'h00f;
rom[411] = 12'h00f;
rom[412] = 12'h00f;
rom[413] = 12'h00f;
rom[414] = 12'h000;
rom[415] = 12'h000;
rom[416] = 12'h000;
rom[417] = 12'h000;
rom[418] = 12'h00f;
rom[419] = 12'h00f;
rom[420] = 12'h00f;
rom[421] = 12'h00f;
rom[422] = 12'h00f;
rom[423] = 12'h00f;
rom[424] = 12'h000;
rom[425] = 12'h000;
rom[426] = 12'h000;
rom[427] = 12'h000;
rom[428] = 12'h000;
rom[429] = 12'h000;
rom[430] = 12'h000;
rom[431] = 12'h000;
rom[432] = 12'h000;
rom[433] = 12'h000;
rom[434] = 12'h00f;
rom[435] = 12'h00f;
rom[436] = 12'h00f;
rom[437] = 12'h00f;
rom[438] = 12'h00f;
rom[439] = 12'h00f;
rom[440] = 12'h000;
rom[441] = 12'h000;
rom[442] = 12'h000;
rom[443] = 12'h000;
rom[444] = 12'h00f;
rom[445] = 12'h00f;
rom[446] = 12'h00f;
rom[447] = 12'h00f;
rom[448] = 12'h00f;
rom[449] = 12'h00f;
rom[450] = 12'h000;
rom[451] = 12'h000;
rom[452] = 12'h000;
rom[453] = 12'h000;
rom[454] = 12'h000;
rom[455] = 12'h000;
rom[456] = 12'h000;
rom[457] = 12'h000;
rom[458] = 12'h000;
rom[459] = 12'h000;
rom[460] = 12'h00f;
rom[461] = 12'h00f;
rom[462] = 12'h00f;
rom[463] = 12'h00f;
rom[464] = 12'h00f;
rom[465] = 12'h00f;
rom[466] = 12'h000;
rom[467] = 12'h000;
rom[468] = 12'h000;
rom[469] = 12'h000;
rom[470] = 12'h00f;
rom[471] = 12'h00f;
rom[472] = 12'h00f;
rom[473] = 12'h00f;
rom[474] = 12'h000;
rom[475] = 12'h000;
rom[476] = 12'h000;
rom[477] = 12'h000;
rom[478] = 12'h000;
rom[479] = 12'h000;
rom[480] = 12'h000;
rom[481] = 12'h000;
rom[482] = 12'h000;
rom[483] = 12'h000;
rom[484] = 12'h000;
rom[485] = 12'h000;
rom[486] = 12'h000;
rom[487] = 12'h000;
rom[488] = 12'h00f;
rom[489] = 12'h00f;
rom[490] = 12'h00f;
rom[491] = 12'h00f;
rom[492] = 12'h000;
rom[493] = 12'h000;
rom[494] = 12'h000;
rom[495] = 12'h000;
rom[496] = 12'h00f;
rom[497] = 12'h00f;
rom[498] = 12'h00f;
rom[499] = 12'h00f;
rom[500] = 12'h000;
rom[501] = 12'h000;
rom[502] = 12'h000;
rom[503] = 12'h000;
rom[504] = 12'h000;
rom[505] = 12'h000;
rom[506] = 12'h000;
rom[507] = 12'h000;
rom[508] = 12'h000;
rom[509] = 12'h000;
rom[510] = 12'h000;
rom[511] = 12'h000;
rom[512] = 12'h000;
rom[513] = 12'h000;
rom[514] = 12'h00f;
rom[515] = 12'h00f;
rom[516] = 12'h00f;
rom[517] = 12'h00f;
rom[518] = 12'h000;
rom[519] = 12'h000;
rom[520] = 12'h000;
rom[521] = 12'h000;
rom[522] = 12'h00f;
rom[523] = 12'h00f;
rom[524] = 12'h000;
rom[525] = 12'h000;
rom[526] = 12'h00f;
rom[527] = 12'h00f;
rom[528] = 12'h00f;
rom[529] = 12'h00f;
rom[530] = 12'h00f;
rom[531] = 12'h00f;
rom[532] = 12'h00f;
rom[533] = 12'h00f;
rom[534] = 12'h00f;
rom[535] = 12'h00f;
rom[536] = 12'h00f;
rom[537] = 12'h00f;
rom[538] = 12'h00f;
rom[539] = 12'h00f;
rom[540] = 12'h000;
rom[541] = 12'h000;
rom[542] = 12'h00f;
rom[543] = 12'h00f;
rom[544] = 12'h000;
rom[545] = 12'h000;
rom[546] = 12'h000;
rom[547] = 12'h000;
rom[548] = 12'h00f;
rom[549] = 12'h00f;
rom[550] = 12'h000;
rom[551] = 12'h000;
rom[552] = 12'h00f;
rom[553] = 12'h00f;
rom[554] = 12'h00f;
rom[555] = 12'h00f;
rom[556] = 12'h00f;
rom[557] = 12'h00f;
rom[558] = 12'h00f;
rom[559] = 12'h00f;
rom[560] = 12'h00f;
rom[561] = 12'h00f;
rom[562] = 12'h00f;
rom[563] = 12'h00f;
rom[564] = 12'h00f;
rom[565] = 12'h00f;
rom[566] = 12'h000;
rom[567] = 12'h000;
rom[568] = 12'h00f;
rom[569] = 12'h00f;
rom[570] = 12'h000;
rom[571] = 12'h000;
rom[572] = 12'h000;
rom[573] = 12'h000;
rom[574] = 12'h000;
rom[575] = 12'h000;
rom[576] = 12'h00f;
rom[577] = 12'h00f;
rom[578] = 12'h00f;
rom[579] = 12'h00f;
rom[580] = 12'h00f;
rom[581] = 12'h00f;
rom[582] = 12'h00f;
rom[583] = 12'h00f;
rom[584] = 12'h00f;
rom[585] = 12'h00f;
rom[586] = 12'h00f;
rom[587] = 12'h00f;
rom[588] = 12'h00f;
rom[589] = 12'h00f;
rom[590] = 12'h00f;
rom[591] = 12'h00f;
rom[592] = 12'h00f;
rom[593] = 12'h00f;
rom[594] = 12'h000;
rom[595] = 12'h000;
rom[596] = 12'h000;
rom[597] = 12'h000;
rom[598] = 12'h000;
rom[599] = 12'h000;
rom[600] = 12'h000;
rom[601] = 12'h000;
rom[602] = 12'h00f;
rom[603] = 12'h00f;
rom[604] = 12'h00f;
rom[605] = 12'h00f;
rom[606] = 12'h00f;
rom[607] = 12'h00f;
rom[608] = 12'h00f;
rom[609] = 12'h00f;
rom[610] = 12'h00f;
rom[611] = 12'h00f;
rom[612] = 12'h00f;
rom[613] = 12'h00f;
rom[614] = 12'h00f;
rom[615] = 12'h00f;
rom[616] = 12'h00f;
rom[617] = 12'h00f;
rom[618] = 12'h00f;
rom[619] = 12'h00f;
rom[620] = 12'h000;
rom[621] = 12'h000;
rom[622] = 12'h000;
rom[623] = 12'h000;
rom[624] = 12'h000;
rom[625] = 12'h000;
rom[626] = 12'h00f;
rom[627] = 12'h00f;
rom[628] = 12'h000;
rom[629] = 12'h000;
rom[630] = 12'h00f;
rom[631] = 12'h00f;
rom[632] = 12'h00f;
rom[633] = 12'h00f;
rom[634] = 12'h00f;
rom[635] = 12'h00f;
rom[636] = 12'h00f;
rom[637] = 12'h00f;
rom[638] = 12'h00f;
rom[639] = 12'h00f;
rom[640] = 12'h00f;
rom[641] = 12'h00f;
rom[642] = 12'h00f;
rom[643] = 12'h00f;
rom[644] = 12'h000;
rom[645] = 12'h000;
rom[646] = 12'h00f;
rom[647] = 12'h00f;
rom[648] = 12'h000;
rom[649] = 12'h000;
rom[650] = 12'h000;
rom[651] = 12'h000;
rom[652] = 12'h00f;
rom[653] = 12'h00f;
rom[654] = 12'h000;
rom[655] = 12'h000;
rom[656] = 12'h00f;
rom[657] = 12'h00f;
rom[658] = 12'h00f;
rom[659] = 12'h00f;
rom[660] = 12'h00f;
rom[661] = 12'h00f;
rom[662] = 12'h00f;
rom[663] = 12'h00f;
rom[664] = 12'h00f;
rom[665] = 12'h00f;
rom[666] = 12'h00f;
rom[667] = 12'h00f;
rom[668] = 12'h00f;
rom[669] = 12'h00f;
rom[670] = 12'h000;
rom[671] = 12'h000;
rom[672] = 12'h00f;
rom[673] = 12'h00f;
rom[674] = 12'h000;
rom[675] = 12'h000;
rom[676] = 12'h000;
rom[677] = 12'h000;
rom[678] = 12'h00f;
rom[679] = 12'h00f;
rom[680] = 12'h00f;
rom[681] = 12'h00f;
rom[682] = 12'h000;
rom[683] = 12'h000;
rom[684] = 12'h000;
rom[685] = 12'h000;
rom[686] = 12'h000;
rom[687] = 12'h000;
rom[688] = 12'h000;
rom[689] = 12'h000;
rom[690] = 12'h000;
rom[691] = 12'h000;
rom[692] = 12'h000;
rom[693] = 12'h000;
rom[694] = 12'h000;
rom[695] = 12'h000;
rom[696] = 12'h00f;
rom[697] = 12'h00f;
rom[698] = 12'h00f;
rom[699] = 12'h00f;
rom[700] = 12'h000;
rom[701] = 12'h000;
rom[702] = 12'h000;
rom[703] = 12'h000;
rom[704] = 12'h00f;
rom[705] = 12'h00f;
rom[706] = 12'h00f;
rom[707] = 12'h00f;
rom[708] = 12'h000;
rom[709] = 12'h000;
rom[710] = 12'h000;
rom[711] = 12'h000;
rom[712] = 12'h000;
rom[713] = 12'h000;
rom[714] = 12'h000;
rom[715] = 12'h000;
rom[716] = 12'h000;
rom[717] = 12'h000;
rom[718] = 12'h000;
rom[719] = 12'h000;
rom[720] = 12'h000;
rom[721] = 12'h000;
rom[722] = 12'h00f;
rom[723] = 12'h00f;
rom[724] = 12'h00f;
rom[725] = 12'h00f;
rom[726] = 12'h000;
rom[727] = 12'h000;
rom[728] = 12'h000;
rom[729] = 12'h000;
rom[730] = 12'h00f;
rom[731] = 12'h00f;
rom[732] = 12'h00f;
rom[733] = 12'h00f;
rom[734] = 12'h00f;
rom[735] = 12'h00f;
rom[736] = 12'h000;
rom[737] = 12'h000;
rom[738] = 12'h000;
rom[739] = 12'h000;
rom[740] = 12'h000;
rom[741] = 12'h000;
rom[742] = 12'h000;
rom[743] = 12'h000;
rom[744] = 12'h000;
rom[745] = 12'h000;
rom[746] = 12'h00f;
rom[747] = 12'h00f;
rom[748] = 12'h00f;
rom[749] = 12'h00f;
rom[750] = 12'h00f;
rom[751] = 12'h00f;
rom[752] = 12'h000;
rom[753] = 12'h000;
rom[754] = 12'h000;
rom[755] = 12'h000;
rom[756] = 12'h00f;
rom[757] = 12'h00f;
rom[758] = 12'h00f;
rom[759] = 12'h00f;
rom[760] = 12'h00f;
rom[761] = 12'h00f;
rom[762] = 12'h000;
rom[763] = 12'h000;
rom[764] = 12'h000;
rom[765] = 12'h000;
rom[766] = 12'h000;
rom[767] = 12'h000;
rom[768] = 12'h000;
rom[769] = 12'h000;
rom[770] = 12'h000;
rom[771] = 12'h000;
rom[772] = 12'h00f;
rom[773] = 12'h00f;
rom[774] = 12'h00f;
rom[775] = 12'h00f;
rom[776] = 12'h00f;
rom[777] = 12'h00f;
rom[778] = 12'h000;
rom[779] = 12'h000;
rom[780] = 12'h000;
rom[781] = 12'h000;
rom[782] = 12'h00f;
rom[783] = 12'h00f;
rom[784] = 12'h00f;
rom[785] = 12'h00f;
rom[786] = 12'h00f;
rom[787] = 12'h00f;
rom[788] = 12'h000;
rom[789] = 12'h000;
rom[790] = 12'h000;
rom[791] = 12'h000;
rom[792] = 12'h000;
rom[793] = 12'h000;
rom[794] = 12'h000;
rom[795] = 12'h000;
rom[796] = 12'h000;
rom[797] = 12'h000;
rom[798] = 12'h00f;
rom[799] = 12'h00f;
rom[800] = 12'h00f;
rom[801] = 12'h00f;
rom[802] = 12'h00f;
rom[803] = 12'h00f;
rom[804] = 12'h000;
rom[805] = 12'h000;
rom[806] = 12'h000;
rom[807] = 12'h000;
rom[808] = 12'h00f;
rom[809] = 12'h00f;
rom[810] = 12'h00f;
rom[811] = 12'h00f;
rom[812] = 12'h00f;
rom[813] = 12'h00f;
rom[814] = 12'h000;
rom[815] = 12'h000;
rom[816] = 12'h000;
rom[817] = 12'h000;
rom[818] = 12'h000;
rom[819] = 12'h000;
rom[820] = 12'h000;
rom[821] = 12'h000;
rom[822] = 12'h000;
rom[823] = 12'h000;
rom[824] = 12'h00f;
rom[825] = 12'h00f;
rom[826] = 12'h00f;
rom[827] = 12'h00f;
rom[828] = 12'h00f;
rom[829] = 12'h00f;
rom[830] = 12'h000;
rom[831] = 12'h000;
rom[832] = 12'h000;
rom[833] = 12'h000;
rom[834] = 12'h00f;
rom[835] = 12'h00f;
rom[836] = 12'h00f;
rom[837] = 12'h00f;
rom[838] = 12'h00f;
rom[839] = 12'h00f;
rom[840] = 12'h000;
rom[841] = 12'h000;
rom[842] = 12'h000;
rom[843] = 12'h000;
rom[844] = 12'h000;
rom[845] = 12'h000;
rom[846] = 12'h000;
rom[847] = 12'h000;
rom[848] = 12'h000;
rom[849] = 12'h000;
rom[850] = 12'h00f;
rom[851] = 12'h00f;
rom[852] = 12'h00f;
rom[853] = 12'h00f;
rom[854] = 12'h00f;
rom[855] = 12'h00f;
rom[856] = 12'h000;
rom[857] = 12'h000;
rom[858] = 12'h000;
rom[859] = 12'h000;
rom[860] = 12'h00f;
rom[861] = 12'h00f;
rom[862] = 12'h00f;
rom[863] = 12'h00f;
rom[864] = 12'h00f;
rom[865] = 12'h00f;
rom[866] = 12'h000;
rom[867] = 12'h000;
rom[868] = 12'h000;
rom[869] = 12'h000;
rom[870] = 12'h000;
rom[871] = 12'h000;
rom[872] = 12'h000;
rom[873] = 12'h000;
rom[874] = 12'h000;
rom[875] = 12'h000;
rom[876] = 12'h00f;
rom[877] = 12'h00f;
rom[878] = 12'h00f;
rom[879] = 12'h00f;
rom[880] = 12'h00f;
rom[881] = 12'h00f;
rom[882] = 12'h000;
rom[883] = 12'h000;
rom[884] = 12'h000;
rom[885] = 12'h000;
rom[886] = 12'h00f;
rom[887] = 12'h00f;
rom[888] = 12'h00f;
rom[889] = 12'h00f;
rom[890] = 12'h00f;
rom[891] = 12'h00f;
rom[892] = 12'h000;
rom[893] = 12'h000;
rom[894] = 12'h000;
rom[895] = 12'h000;
rom[896] = 12'h000;
rom[897] = 12'h000;
rom[898] = 12'h000;
rom[899] = 12'h000;
rom[900] = 12'h000;
rom[901] = 12'h000;
rom[902] = 12'h00f;
rom[903] = 12'h00f;
rom[904] = 12'h00f;
rom[905] = 12'h00f;
rom[906] = 12'h00f;
rom[907] = 12'h00f;
rom[908] = 12'h000;
rom[909] = 12'h000;
rom[910] = 12'h000;
rom[911] = 12'h000;
rom[912] = 12'h00f;
rom[913] = 12'h00f;
rom[914] = 12'h00f;
rom[915] = 12'h00f;
rom[916] = 12'h00f;
rom[917] = 12'h00f;
rom[918] = 12'h000;
rom[919] = 12'h000;
rom[920] = 12'h000;
rom[921] = 12'h000;
rom[922] = 12'h000;
rom[923] = 12'h000;
rom[924] = 12'h000;
rom[925] = 12'h000;
rom[926] = 12'h000;
rom[927] = 12'h000;
rom[928] = 12'h00f;
rom[929] = 12'h00f;
rom[930] = 12'h00f;
rom[931] = 12'h00f;
rom[932] = 12'h00f;
rom[933] = 12'h00f;
rom[934] = 12'h000;
rom[935] = 12'h000;
rom[936] = 12'h000;
rom[937] = 12'h000;
rom[938] = 12'h00f;
rom[939] = 12'h00f;
rom[940] = 12'h00f;
rom[941] = 12'h00f;
rom[942] = 12'h00f;
rom[943] = 12'h00f;
rom[944] = 12'h000;
rom[945] = 12'h000;
rom[946] = 12'h000;
rom[947] = 12'h000;
rom[948] = 12'h000;
rom[949] = 12'h000;
rom[950] = 12'h000;
rom[951] = 12'h000;
rom[952] = 12'h000;
rom[953] = 12'h000;
rom[954] = 12'h00f;
rom[955] = 12'h00f;
rom[956] = 12'h00f;
rom[957] = 12'h00f;
rom[958] = 12'h00f;
rom[959] = 12'h00f;
rom[960] = 12'h000;
rom[961] = 12'h000;
rom[962] = 12'h000;
rom[963] = 12'h000;
rom[964] = 12'h00f;
rom[965] = 12'h00f;
rom[966] = 12'h00f;
rom[967] = 12'h00f;
rom[968] = 12'h00f;
rom[969] = 12'h00f;
rom[970] = 12'h000;
rom[971] = 12'h000;
rom[972] = 12'h000;
rom[973] = 12'h000;
rom[974] = 12'h000;
rom[975] = 12'h000;
rom[976] = 12'h000;
rom[977] = 12'h000;
rom[978] = 12'h000;
rom[979] = 12'h000;
rom[980] = 12'h00f;
rom[981] = 12'h00f;
rom[982] = 12'h00f;
rom[983] = 12'h00f;
rom[984] = 12'h00f;
rom[985] = 12'h00f;
rom[986] = 12'h000;
rom[987] = 12'h000;
rom[988] = 12'h000;
rom[989] = 12'h000;
rom[990] = 12'h00f;
rom[991] = 12'h00f;
rom[992] = 12'h00f;
rom[993] = 12'h00f;
rom[994] = 12'h000;
rom[995] = 12'h000;
rom[996] = 12'h00f;
rom[997] = 12'h00f;
rom[998] = 12'h00f;
rom[999] = 12'h00f;
rom[1000] = 12'h00f;
rom[1001] = 12'h00f;
rom[1002] = 12'h00f;
rom[1003] = 12'h00f;
rom[1004] = 12'h00f;
rom[1005] = 12'h00f;
rom[1006] = 12'h000;
rom[1007] = 12'h000;
rom[1008] = 12'h00f;
rom[1009] = 12'h00f;
rom[1010] = 12'h00f;
rom[1011] = 12'h00f;
rom[1012] = 12'h000;
rom[1013] = 12'h000;
rom[1014] = 12'h000;
rom[1015] = 12'h000;
rom[1016] = 12'h00f;
rom[1017] = 12'h00f;
rom[1018] = 12'h00f;
rom[1019] = 12'h00f;
rom[1020] = 12'h000;
rom[1021] = 12'h000;
rom[1022] = 12'h00f;
rom[1023] = 12'h00f;
rom[1024] = 12'h00f;
rom[1025] = 12'h00f;
rom[1026] = 12'h00f;
rom[1027] = 12'h00f;
rom[1028] = 12'h00f;
rom[1029] = 12'h00f;
rom[1030] = 12'h00f;
rom[1031] = 12'h00f;
rom[1032] = 12'h000;
rom[1033] = 12'h000;
rom[1034] = 12'h00f;
rom[1035] = 12'h00f;
rom[1036] = 12'h00f;
rom[1037] = 12'h00f;
rom[1038] = 12'h000;
rom[1039] = 12'h000;
rom[1040] = 12'h000;
rom[1041] = 12'h000;
rom[1042] = 12'h00f;
rom[1043] = 12'h00f;
rom[1044] = 12'h000;
rom[1045] = 12'h000;
rom[1046] = 12'h00f;
rom[1047] = 12'h00f;
rom[1048] = 12'h00f;
rom[1049] = 12'h00f;
rom[1050] = 12'h00f;
rom[1051] = 12'h00f;
rom[1052] = 12'h00f;
rom[1053] = 12'h00f;
rom[1054] = 12'h00f;
rom[1055] = 12'h00f;
rom[1056] = 12'h00f;
rom[1057] = 12'h00f;
rom[1058] = 12'h00f;
rom[1059] = 12'h00f;
rom[1060] = 12'h000;
rom[1061] = 12'h000;
rom[1062] = 12'h00f;
rom[1063] = 12'h00f;
rom[1064] = 12'h000;
rom[1065] = 12'h000;
rom[1066] = 12'h000;
rom[1067] = 12'h000;
rom[1068] = 12'h00f;
rom[1069] = 12'h00f;
rom[1070] = 12'h000;
rom[1071] = 12'h000;
rom[1072] = 12'h00f;
rom[1073] = 12'h00f;
rom[1074] = 12'h00f;
rom[1075] = 12'h00f;
rom[1076] = 12'h00f;
rom[1077] = 12'h00f;
rom[1078] = 12'h00f;
rom[1079] = 12'h00f;
rom[1080] = 12'h00f;
rom[1081] = 12'h00f;
rom[1082] = 12'h00f;
rom[1083] = 12'h00f;
rom[1084] = 12'h00f;
rom[1085] = 12'h00f;
rom[1086] = 12'h000;
rom[1087] = 12'h000;
rom[1088] = 12'h00f;
rom[1089] = 12'h00f;
rom[1090] = 12'h000;
rom[1091] = 12'h000;
rom[1092] = 12'h000;
rom[1093] = 12'h000;
rom[1094] = 12'h000;
rom[1095] = 12'h000;
rom[1096] = 12'h00f;
rom[1097] = 12'h00f;
rom[1098] = 12'h00f;
rom[1099] = 12'h00f;
rom[1100] = 12'h00f;
rom[1101] = 12'h00f;
rom[1102] = 12'h00f;
rom[1103] = 12'h00f;
rom[1104] = 12'h00f;
rom[1105] = 12'h00f;
rom[1106] = 12'h00f;
rom[1107] = 12'h00f;
rom[1108] = 12'h00f;
rom[1109] = 12'h00f;
rom[1110] = 12'h00f;
rom[1111] = 12'h00f;
rom[1112] = 12'h00f;
rom[1113] = 12'h00f;
rom[1114] = 12'h000;
rom[1115] = 12'h000;
rom[1116] = 12'h000;
rom[1117] = 12'h000;
rom[1118] = 12'h000;
rom[1119] = 12'h000;
rom[1120] = 12'h000;
rom[1121] = 12'h000;
rom[1122] = 12'h00f;
rom[1123] = 12'h00f;
rom[1124] = 12'h00f;
rom[1125] = 12'h00f;
rom[1126] = 12'h00f;
rom[1127] = 12'h00f;
rom[1128] = 12'h00f;
rom[1129] = 12'h00f;
rom[1130] = 12'h00f;
rom[1131] = 12'h00f;
rom[1132] = 12'h00f;
rom[1133] = 12'h00f;
rom[1134] = 12'h00f;
rom[1135] = 12'h00f;
rom[1136] = 12'h00f;
rom[1137] = 12'h00f;
rom[1138] = 12'h00f;
rom[1139] = 12'h00f;
rom[1140] = 12'h000;
rom[1141] = 12'h000;
rom[1142] = 12'h000;
rom[1143] = 12'h000;
rom[1144] = 12'h000;
rom[1145] = 12'h000;
rom[1146] = 12'h000;
rom[1147] = 12'h000;
rom[1148] = 12'h000;
rom[1149] = 12'h000;
rom[1150] = 12'h000;
rom[1151] = 12'h000;
rom[1152] = 12'h000;
rom[1153] = 12'h000;
rom[1154] = 12'h000;
rom[1155] = 12'h000;
rom[1156] = 12'h000;
rom[1157] = 12'h000;
rom[1158] = 12'h000;
rom[1159] = 12'h000;
rom[1160] = 12'h000;
rom[1161] = 12'h000;
rom[1162] = 12'h000;
rom[1163] = 12'h000;
rom[1164] = 12'h000;
rom[1165] = 12'h000;
rom[1166] = 12'h000;
rom[1167] = 12'h000;
rom[1168] = 12'h000;
rom[1169] = 12'h000;
rom[1170] = 12'h000;
rom[1171] = 12'h000;
rom[1172] = 12'h000;
rom[1173] = 12'h000;
rom[1174] = 12'h000;
rom[1175] = 12'h000;
rom[1176] = 12'h000;
rom[1177] = 12'h000;
rom[1178] = 12'h000;
rom[1179] = 12'h000;
rom[1180] = 12'h000;
rom[1181] = 12'h000;
rom[1182] = 12'h000;
rom[1183] = 12'h000;
rom[1184] = 12'h000;
rom[1185] = 12'h000;
rom[1186] = 12'h000;
rom[1187] = 12'h000;
rom[1188] = 12'h000;
rom[1189] = 12'h000;
rom[1190] = 12'h000;
rom[1191] = 12'h000;
rom[1192] = 12'h000;
rom[1193] = 12'h000;
rom[1194] = 12'h000;
rom[1195] = 12'h000;

  end
  endmodule

    module dash_rom (                       //девять
  input  wire    [13:0]     addr,
  output wire    [11:0]     word
);

  logic [11:0] rom [(25 * 25)];

  assign word = rom[addr];

  initial begin
rom[0] = 12'h000;
rom[1] = 12'h000;
rom[2] = 12'h000;
rom[3] = 12'h000;
rom[4] = 12'h000;
rom[5] = 12'h000;
rom[6] = 12'h000;
rom[7] = 12'h000;
rom[8] = 12'h000;
rom[9] = 12'h000;
rom[10] = 12'h000;
rom[11] = 12'h000;
rom[12] = 12'h000;
rom[13] = 12'h000;
rom[14] = 12'h000;
rom[15] = 12'h000;
rom[16] = 12'h000;
rom[17] = 12'h000;
rom[18] = 12'h000;
rom[19] = 12'h000;
rom[20] = 12'h000;
rom[21] = 12'h000;
rom[22] = 12'h000;
rom[23] = 12'h000;
rom[24] = 12'h000;
rom[25] = 12'h000;
rom[26] = 12'h000;
rom[27] = 12'h000;
rom[28] = 12'h000;
rom[29] = 12'h000;
rom[30] = 12'h000;
rom[31] = 12'h000;
rom[32] = 12'h000;
rom[33] = 12'h000;
rom[34] = 12'h000;
rom[35] = 12'h000;
rom[36] = 12'h000;
rom[37] = 12'h000;
rom[38] = 12'h000;
rom[39] = 12'h000;
rom[40] = 12'h000;
rom[41] = 12'h000;
rom[42] = 12'h000;
rom[43] = 12'h000;
rom[44] = 12'h000;
rom[45] = 12'h000;
rom[46] = 12'h000;
rom[47] = 12'h000;
rom[48] = 12'h000;
rom[49] = 12'h000;
rom[50] = 12'h000;
rom[51] = 12'h000;
rom[52] = 12'h000;
rom[53] = 12'h000;
rom[54] = 12'h000;
rom[55] = 12'h000;
rom[56] = 12'h00f;
rom[57] = 12'h00f;
rom[58] = 12'h00f;
rom[59] = 12'h00f;
rom[60] = 12'h00f;
rom[61] = 12'h00f;
rom[62] = 12'h00f;
rom[63] = 12'h00f;
rom[64] = 12'h00f;
rom[65] = 12'h00f;
rom[66] = 12'h00f;
rom[67] = 12'h00f;
rom[68] = 12'h00f;
rom[69] = 12'h00f;
rom[70] = 12'h00f;
rom[71] = 12'h00f;
rom[72] = 12'h00f;
rom[73] = 12'h00f;
rom[74] = 12'h000;
rom[75] = 12'h000;
rom[76] = 12'h000;
rom[77] = 12'h000;
rom[78] = 12'h000;
rom[79] = 12'h000;
rom[80] = 12'h000;
rom[81] = 12'h000;
rom[82] = 12'h00f;
rom[83] = 12'h00f;
rom[84] = 12'h00f;
rom[85] = 12'h00f;
rom[86] = 12'h00f;
rom[87] = 12'h00f;
rom[88] = 12'h00f;
rom[89] = 12'h00f;
rom[90] = 12'h00f;
rom[91] = 12'h00f;
rom[92] = 12'h00f;
rom[93] = 12'h00f;
rom[94] = 12'h00f;
rom[95] = 12'h00f;
rom[96] = 12'h00f;
rom[97] = 12'h00f;
rom[98] = 12'h00f;
rom[99] = 12'h00f;
rom[100] = 12'h000;
rom[101] = 12'h000;
rom[102] = 12'h000;
rom[103] = 12'h000;
rom[104] = 12'h000;
rom[105] = 12'h000;
rom[106] = 12'h00f;
rom[107] = 12'h00f;
rom[108] = 12'h000;
rom[109] = 12'h000;
rom[110] = 12'h00f;
rom[111] = 12'h00f;
rom[112] = 12'h00f;
rom[113] = 12'h00f;
rom[114] = 12'h00f;
rom[115] = 12'h00f;
rom[116] = 12'h00f;
rom[117] = 12'h00f;
rom[118] = 12'h00f;
rom[119] = 12'h00f;
rom[120] = 12'h00f;
rom[121] = 12'h00f;
rom[122] = 12'h00f;
rom[123] = 12'h00f;
rom[124] = 12'h000;
rom[125] = 12'h000;
rom[126] = 12'h00f;
rom[127] = 12'h00f;
rom[128] = 12'h000;
rom[129] = 12'h000;
rom[130] = 12'h000;
rom[131] = 12'h000;
rom[132] = 12'h00f;
rom[133] = 12'h00f;
rom[134] = 12'h000;
rom[135] = 12'h000;
rom[136] = 12'h00f;
rom[137] = 12'h00f;
rom[138] = 12'h00f;
rom[139] = 12'h00f;
rom[140] = 12'h00f;
rom[141] = 12'h00f;
rom[142] = 12'h00f;
rom[143] = 12'h00f;
rom[144] = 12'h00f;
rom[145] = 12'h00f;
rom[146] = 12'h00f;
rom[147] = 12'h00f;
rom[148] = 12'h00f;
rom[149] = 12'h00f;
rom[150] = 12'h000;
rom[151] = 12'h000;
rom[152] = 12'h00f;
rom[153] = 12'h00f;
rom[154] = 12'h000;
rom[155] = 12'h000;
rom[156] = 12'h000;
rom[157] = 12'h000;
rom[158] = 12'h00f;
rom[159] = 12'h00f;
rom[160] = 12'h00f;
rom[161] = 12'h00f;
rom[162] = 12'h000;
rom[163] = 12'h000;
rom[164] = 12'h00f;
rom[165] = 12'h00f;
rom[166] = 12'h00f;
rom[167] = 12'h00f;
rom[168] = 12'h00f;
rom[169] = 12'h00f;
rom[170] = 12'h00f;
rom[171] = 12'h00f;
rom[172] = 12'h00f;
rom[173] = 12'h00f;
rom[174] = 12'h000;
rom[175] = 12'h000;
rom[176] = 12'h00f;
rom[177] = 12'h00f;
rom[178] = 12'h00f;
rom[179] = 12'h00f;
rom[180] = 12'h000;
rom[181] = 12'h000;
rom[182] = 12'h000;
rom[183] = 12'h000;
rom[184] = 12'h00f;
rom[185] = 12'h00f;
rom[186] = 12'h00f;
rom[187] = 12'h00f;
rom[188] = 12'h000;
rom[189] = 12'h000;
rom[190] = 12'h00f;
rom[191] = 12'h00f;
rom[192] = 12'h00f;
rom[193] = 12'h00f;
rom[194] = 12'h00f;
rom[195] = 12'h00f;
rom[196] = 12'h00f;
rom[197] = 12'h00f;
rom[198] = 12'h00f;
rom[199] = 12'h00f;
rom[200] = 12'h000;
rom[201] = 12'h000;
rom[202] = 12'h00f;
rom[203] = 12'h00f;
rom[204] = 12'h00f;
rom[205] = 12'h00f;
rom[206] = 12'h000;
rom[207] = 12'h000;
rom[208] = 12'h000;
rom[209] = 12'h000;
rom[210] = 12'h00f;
rom[211] = 12'h00f;
rom[212] = 12'h00f;
rom[213] = 12'h00f;
rom[214] = 12'h00f;
rom[215] = 12'h00f;
rom[216] = 12'h000;
rom[217] = 12'h000;
rom[218] = 12'h000;
rom[219] = 12'h000;
rom[220] = 12'h000;
rom[221] = 12'h000;
rom[222] = 12'h000;
rom[223] = 12'h000;
rom[224] = 12'h000;
rom[225] = 12'h000;
rom[226] = 12'h00f;
rom[227] = 12'h00f;
rom[228] = 12'h00f;
rom[229] = 12'h00f;
rom[230] = 12'h00f;
rom[231] = 12'h00f;
rom[232] = 12'h000;
rom[233] = 12'h000;
rom[234] = 12'h000;
rom[235] = 12'h000;
rom[236] = 12'h00f;
rom[237] = 12'h00f;
rom[238] = 12'h00f;
rom[239] = 12'h00f;
rom[240] = 12'h00f;
rom[241] = 12'h00f;
rom[242] = 12'h000;
rom[243] = 12'h000;
rom[244] = 12'h000;
rom[245] = 12'h000;
rom[246] = 12'h000;
rom[247] = 12'h000;
rom[248] = 12'h000;
rom[249] = 12'h000;
rom[250] = 12'h000;
rom[251] = 12'h000;
rom[252] = 12'h00f;
rom[253] = 12'h00f;
rom[254] = 12'h00f;
rom[255] = 12'h00f;
rom[256] = 12'h00f;
rom[257] = 12'h00f;
rom[258] = 12'h000;
rom[259] = 12'h000;
rom[260] = 12'h000;
rom[261] = 12'h000;
rom[262] = 12'h00f;
rom[263] = 12'h00f;
rom[264] = 12'h00f;
rom[265] = 12'h00f;
rom[266] = 12'h00f;
rom[267] = 12'h00f;
rom[268] = 12'h000;
rom[269] = 12'h000;
rom[270] = 12'h000;
rom[271] = 12'h000;
rom[272] = 12'h000;
rom[273] = 12'h000;
rom[274] = 12'h000;
rom[275] = 12'h000;
rom[276] = 12'h000;
rom[277] = 12'h000;
rom[278] = 12'h00f;
rom[279] = 12'h00f;
rom[280] = 12'h00f;
rom[281] = 12'h00f;
rom[282] = 12'h00f;
rom[283] = 12'h00f;
rom[284] = 12'h000;
rom[285] = 12'h000;
rom[286] = 12'h000;
rom[287] = 12'h000;
rom[288] = 12'h00f;
rom[289] = 12'h00f;
rom[290] = 12'h00f;
rom[291] = 12'h00f;
rom[292] = 12'h00f;
rom[293] = 12'h00f;
rom[294] = 12'h000;
rom[295] = 12'h000;
rom[296] = 12'h000;
rom[297] = 12'h000;
rom[298] = 12'h000;
rom[299] = 12'h000;
rom[300] = 12'h000;
rom[301] = 12'h000;
rom[302] = 12'h000;
rom[303] = 12'h000;
rom[304] = 12'h00f;
rom[305] = 12'h00f;
rom[306] = 12'h00f;
rom[307] = 12'h00f;
rom[308] = 12'h00f;
rom[309] = 12'h00f;
rom[310] = 12'h000;
rom[311] = 12'h000;
rom[312] = 12'h000;
rom[313] = 12'h000;
rom[314] = 12'h00f;
rom[315] = 12'h00f;
rom[316] = 12'h00f;
rom[317] = 12'h00f;
rom[318] = 12'h00f;
rom[319] = 12'h00f;
rom[320] = 12'h000;
rom[321] = 12'h000;
rom[322] = 12'h000;
rom[323] = 12'h000;
rom[324] = 12'h000;
rom[325] = 12'h000;
rom[326] = 12'h000;
rom[327] = 12'h000;
rom[328] = 12'h000;
rom[329] = 12'h000;
rom[330] = 12'h00f;
rom[331] = 12'h00f;
rom[332] = 12'h00f;
rom[333] = 12'h00f;
rom[334] = 12'h00f;
rom[335] = 12'h00f;
rom[336] = 12'h000;
rom[337] = 12'h000;
rom[338] = 12'h000;
rom[339] = 12'h000;
rom[340] = 12'h00f;
rom[341] = 12'h00f;
rom[342] = 12'h00f;
rom[343] = 12'h00f;
rom[344] = 12'h00f;
rom[345] = 12'h00f;
rom[346] = 12'h000;
rom[347] = 12'h000;
rom[348] = 12'h000;
rom[349] = 12'h000;
rom[350] = 12'h000;
rom[351] = 12'h000;
rom[352] = 12'h000;
rom[353] = 12'h000;
rom[354] = 12'h000;
rom[355] = 12'h000;
rom[356] = 12'h00f;
rom[357] = 12'h00f;
rom[358] = 12'h00f;
rom[359] = 12'h00f;
rom[360] = 12'h00f;
rom[361] = 12'h00f;
rom[362] = 12'h000;
rom[363] = 12'h000;
rom[364] = 12'h000;
rom[365] = 12'h000;
rom[366] = 12'h00f;
rom[367] = 12'h00f;
rom[368] = 12'h00f;
rom[369] = 12'h00f;
rom[370] = 12'h00f;
rom[371] = 12'h00f;
rom[372] = 12'h000;
rom[373] = 12'h000;
rom[374] = 12'h000;
rom[375] = 12'h000;
rom[376] = 12'h000;
rom[377] = 12'h000;
rom[378] = 12'h000;
rom[379] = 12'h000;
rom[380] = 12'h000;
rom[381] = 12'h000;
rom[382] = 12'h00f;
rom[383] = 12'h00f;
rom[384] = 12'h00f;
rom[385] = 12'h00f;
rom[386] = 12'h00f;
rom[387] = 12'h00f;
rom[388] = 12'h000;
rom[389] = 12'h000;
rom[390] = 12'h000;
rom[391] = 12'h000;
rom[392] = 12'h00f;
rom[393] = 12'h00f;
rom[394] = 12'h00f;
rom[395] = 12'h00f;
rom[396] = 12'h00f;
rom[397] = 12'h00f;
rom[398] = 12'h000;
rom[399] = 12'h000;
rom[400] = 12'h000;
rom[401] = 12'h000;
rom[402] = 12'h000;
rom[403] = 12'h000;
rom[404] = 12'h000;
rom[405] = 12'h000;
rom[406] = 12'h000;
rom[407] = 12'h000;
rom[408] = 12'h00f;
rom[409] = 12'h00f;
rom[410] = 12'h00f;
rom[411] = 12'h00f;
rom[412] = 12'h00f;
rom[413] = 12'h00f;
rom[414] = 12'h000;
rom[415] = 12'h000;
rom[416] = 12'h000;
rom[417] = 12'h000;
rom[418] = 12'h00f;
rom[419] = 12'h00f;
rom[420] = 12'h00f;
rom[421] = 12'h00f;
rom[422] = 12'h00f;
rom[423] = 12'h00f;
rom[424] = 12'h000;
rom[425] = 12'h000;
rom[426] = 12'h000;
rom[427] = 12'h000;
rom[428] = 12'h000;
rom[429] = 12'h000;
rom[430] = 12'h000;
rom[431] = 12'h000;
rom[432] = 12'h000;
rom[433] = 12'h000;
rom[434] = 12'h00f;
rom[435] = 12'h00f;
rom[436] = 12'h00f;
rom[437] = 12'h00f;
rom[438] = 12'h00f;
rom[439] = 12'h00f;
rom[440] = 12'h000;
rom[441] = 12'h000;
rom[442] = 12'h000;
rom[443] = 12'h000;
rom[444] = 12'h00f;
rom[445] = 12'h00f;
rom[446] = 12'h00f;
rom[447] = 12'h00f;
rom[448] = 12'h00f;
rom[449] = 12'h00f;
rom[450] = 12'h000;
rom[451] = 12'h000;
rom[452] = 12'h000;
rom[453] = 12'h000;
rom[454] = 12'h000;
rom[455] = 12'h000;
rom[456] = 12'h000;
rom[457] = 12'h000;
rom[458] = 12'h000;
rom[459] = 12'h000;
rom[460] = 12'h00f;
rom[461] = 12'h00f;
rom[462] = 12'h00f;
rom[463] = 12'h00f;
rom[464] = 12'h00f;
rom[465] = 12'h00f;
rom[466] = 12'h000;
rom[467] = 12'h000;
rom[468] = 12'h000;
rom[469] = 12'h000;
rom[470] = 12'h00f;
rom[471] = 12'h00f;
rom[472] = 12'h00f;
rom[473] = 12'h00f;
rom[474] = 12'h000;
rom[475] = 12'h000;
rom[476] = 12'h000;
rom[477] = 12'h000;
rom[478] = 12'h000;
rom[479] = 12'h000;
rom[480] = 12'h000;
rom[481] = 12'h000;
rom[482] = 12'h000;
rom[483] = 12'h000;
rom[484] = 12'h000;
rom[485] = 12'h000;
rom[486] = 12'h000;
rom[487] = 12'h000;
rom[488] = 12'h00f;
rom[489] = 12'h00f;
rom[490] = 12'h00f;
rom[491] = 12'h00f;
rom[492] = 12'h000;
rom[493] = 12'h000;
rom[494] = 12'h000;
rom[495] = 12'h000;
rom[496] = 12'h00f;
rom[497] = 12'h00f;
rom[498] = 12'h00f;
rom[499] = 12'h00f;
rom[500] = 12'h000;
rom[501] = 12'h000;
rom[502] = 12'h000;
rom[503] = 12'h000;
rom[504] = 12'h000;
rom[505] = 12'h000;
rom[506] = 12'h000;
rom[507] = 12'h000;
rom[508] = 12'h000;
rom[509] = 12'h000;
rom[510] = 12'h000;
rom[511] = 12'h000;
rom[512] = 12'h000;
rom[513] = 12'h000;
rom[514] = 12'h00f;
rom[515] = 12'h00f;
rom[516] = 12'h00f;
rom[517] = 12'h00f;
rom[518] = 12'h000;
rom[519] = 12'h000;
rom[520] = 12'h000;
rom[521] = 12'h000;
rom[522] = 12'h00f;
rom[523] = 12'h00f;
rom[524] = 12'h000;
rom[525] = 12'h000;
rom[526] = 12'h00f;
rom[527] = 12'h00f;
rom[528] = 12'h00f;
rom[529] = 12'h00f;
rom[530] = 12'h00f;
rom[531] = 12'h00f;
rom[532] = 12'h00f;
rom[533] = 12'h00f;
rom[534] = 12'h00f;
rom[535] = 12'h00f;
rom[536] = 12'h00f;
rom[537] = 12'h00f;
rom[538] = 12'h00f;
rom[539] = 12'h00f;
rom[540] = 12'h000;
rom[541] = 12'h000;
rom[542] = 12'h00f;
rom[543] = 12'h00f;
rom[544] = 12'h000;
rom[545] = 12'h000;
rom[546] = 12'h000;
rom[547] = 12'h000;
rom[548] = 12'h00f;
rom[549] = 12'h00f;
rom[550] = 12'h000;
rom[551] = 12'h000;
rom[552] = 12'h00f;
rom[553] = 12'h00f;
rom[554] = 12'h00f;
rom[555] = 12'h00f;
rom[556] = 12'h00f;
rom[557] = 12'h00f;
rom[558] = 12'h00f;
rom[559] = 12'h00f;
rom[560] = 12'h00f;
rom[561] = 12'h00f;
rom[562] = 12'h00f;
rom[563] = 12'h00f;
rom[564] = 12'h00f;
rom[565] = 12'h00f;
rom[566] = 12'h000;
rom[567] = 12'h000;
rom[568] = 12'h00f;
rom[569] = 12'h00f;
rom[570] = 12'h000;
rom[571] = 12'h000;
rom[572] = 12'h000;
rom[573] = 12'h000;
rom[574] = 12'h000;
rom[575] = 12'h000;
rom[576] = 12'h00f;
rom[577] = 12'h00f;
rom[578] = 12'h00f;
rom[579] = 12'h00f;
rom[580] = 12'h00f;
rom[581] = 12'h00f;
rom[582] = 12'h00f;
rom[583] = 12'h00f;
rom[584] = 12'h00f;
rom[585] = 12'h00f;
rom[586] = 12'h00f;
rom[587] = 12'h00f;
rom[588] = 12'h00f;
rom[589] = 12'h00f;
rom[590] = 12'h00f;
rom[591] = 12'h00f;
rom[592] = 12'h00f;
rom[593] = 12'h00f;
rom[594] = 12'h000;
rom[595] = 12'h000;
rom[596] = 12'h000;
rom[597] = 12'h000;
rom[598] = 12'h000;
rom[599] = 12'h000;
rom[600] = 12'h000;
rom[601] = 12'h000;
rom[602] = 12'h00f;
rom[603] = 12'h00f;
rom[604] = 12'h00f;
rom[605] = 12'h00f;
rom[606] = 12'h00f;
rom[607] = 12'h00f;
rom[608] = 12'h00f;
rom[609] = 12'h00f;
rom[610] = 12'h00f;
rom[611] = 12'h00f;
rom[612] = 12'h00f;
rom[613] = 12'h00f;
rom[614] = 12'h00f;
rom[615] = 12'h00f;
rom[616] = 12'h00f;
rom[617] = 12'h00f;
rom[618] = 12'h00f;
rom[619] = 12'h00f;
rom[620] = 12'h000;
rom[621] = 12'h000;
rom[622] = 12'h000;
rom[623] = 12'h000;
rom[624] = 12'h000;
rom[625] = 12'h000;
rom[626] = 12'h007;
rom[627] = 12'h007;
rom[628] = 12'h000;
rom[629] = 12'h000;
rom[630] = 12'h00f;
rom[631] = 12'h00f;
rom[632] = 12'h00f;
rom[633] = 12'h00f;
rom[634] = 12'h00f;
rom[635] = 12'h00f;
rom[636] = 12'h00f;
rom[637] = 12'h00f;
rom[638] = 12'h00f;
rom[639] = 12'h00f;
rom[640] = 12'h00f;
rom[641] = 12'h00f;
rom[642] = 12'h00f;
rom[643] = 12'h00f;
rom[644] = 12'h000;
rom[645] = 12'h000;
rom[646] = 12'h00f;
rom[647] = 12'h00f;
rom[648] = 12'h000;
rom[649] = 12'h000;
rom[650] = 12'h000;
rom[651] = 12'h000;
rom[652] = 12'h007;
rom[653] = 12'h007;
rom[654] = 12'h000;
rom[655] = 12'h000;
rom[656] = 12'h00f;
rom[657] = 12'h00f;
rom[658] = 12'h00f;
rom[659] = 12'h00f;
rom[660] = 12'h00f;
rom[661] = 12'h00f;
rom[662] = 12'h00f;
rom[663] = 12'h00f;
rom[664] = 12'h00f;
rom[665] = 12'h00f;
rom[666] = 12'h00f;
rom[667] = 12'h00f;
rom[668] = 12'h00f;
rom[669] = 12'h00f;
rom[670] = 12'h000;
rom[671] = 12'h000;
rom[672] = 12'h00f;
rom[673] = 12'h00f;
rom[674] = 12'h000;
rom[675] = 12'h000;
rom[676] = 12'h000;
rom[677] = 12'h000;
rom[678] = 12'h000;
rom[679] = 12'h000;
rom[680] = 12'h007;
rom[681] = 12'h007;
rom[682] = 12'h000;
rom[683] = 12'h000;
rom[684] = 12'h000;
rom[685] = 12'h000;
rom[686] = 12'h000;
rom[687] = 12'h000;
rom[688] = 12'h000;
rom[689] = 12'h000;
rom[690] = 12'h000;
rom[691] = 12'h000;
rom[692] = 12'h000;
rom[693] = 12'h000;
rom[694] = 12'h000;
rom[695] = 12'h000;
rom[696] = 12'h00f;
rom[697] = 12'h00f;
rom[698] = 12'h00f;
rom[699] = 12'h00f;
rom[700] = 12'h000;
rom[701] = 12'h000;
rom[702] = 12'h000;
rom[703] = 12'h000;
rom[704] = 12'h000;
rom[705] = 12'h000;
rom[706] = 12'h007;
rom[707] = 12'h007;
rom[708] = 12'h000;
rom[709] = 12'h000;
rom[710] = 12'h000;
rom[711] = 12'h000;
rom[712] = 12'h000;
rom[713] = 12'h000;
rom[714] = 12'h000;
rom[715] = 12'h000;
rom[716] = 12'h000;
rom[717] = 12'h000;
rom[718] = 12'h000;
rom[719] = 12'h000;
rom[720] = 12'h000;
rom[721] = 12'h000;
rom[722] = 12'h00f;
rom[723] = 12'h00f;
rom[724] = 12'h00f;
rom[725] = 12'h00f;
rom[726] = 12'h000;
rom[727] = 12'h000;
rom[728] = 12'h000;
rom[729] = 12'h000;
rom[730] = 12'h007;
rom[731] = 12'h007;
rom[732] = 12'h000;
rom[733] = 12'h000;
rom[734] = 12'h007;
rom[735] = 12'h007;
rom[736] = 12'h000;
rom[737] = 12'h000;
rom[738] = 12'h000;
rom[739] = 12'h000;
rom[740] = 12'h000;
rom[741] = 12'h000;
rom[742] = 12'h000;
rom[743] = 12'h000;
rom[744] = 12'h000;
rom[745] = 12'h000;
rom[746] = 12'h00f;
rom[747] = 12'h00f;
rom[748] = 12'h00f;
rom[749] = 12'h00f;
rom[750] = 12'h00f;
rom[751] = 12'h00f;
rom[752] = 12'h000;
rom[753] = 12'h000;
rom[754] = 12'h000;
rom[755] = 12'h000;
rom[756] = 12'h007;
rom[757] = 12'h007;
rom[758] = 12'h000;
rom[759] = 12'h000;
rom[760] = 12'h007;
rom[761] = 12'h007;
rom[762] = 12'h000;
rom[763] = 12'h000;
rom[764] = 12'h000;
rom[765] = 12'h000;
rom[766] = 12'h000;
rom[767] = 12'h000;
rom[768] = 12'h000;
rom[769] = 12'h000;
rom[770] = 12'h000;
rom[771] = 12'h000;
rom[772] = 12'h00f;
rom[773] = 12'h00f;
rom[774] = 12'h00f;
rom[775] = 12'h00f;
rom[776] = 12'h00f;
rom[777] = 12'h00f;
rom[778] = 12'h000;
rom[779] = 12'h000;
rom[780] = 12'h000;
rom[781] = 12'h000;
rom[782] = 12'h000;
rom[783] = 12'h000;
rom[784] = 12'h007;
rom[785] = 12'h007;
rom[786] = 12'h000;
rom[787] = 12'h000;
rom[788] = 12'h000;
rom[789] = 12'h000;
rom[790] = 12'h000;
rom[791] = 12'h000;
rom[792] = 12'h000;
rom[793] = 12'h000;
rom[794] = 12'h000;
rom[795] = 12'h000;
rom[796] = 12'h000;
rom[797] = 12'h000;
rom[798] = 12'h00f;
rom[799] = 12'h00f;
rom[800] = 12'h00f;
rom[801] = 12'h00f;
rom[802] = 12'h00f;
rom[803] = 12'h00f;
rom[804] = 12'h000;
rom[805] = 12'h000;
rom[806] = 12'h000;
rom[807] = 12'h000;
rom[808] = 12'h000;
rom[809] = 12'h000;
rom[810] = 12'h007;
rom[811] = 12'h007;
rom[812] = 12'h000;
rom[813] = 12'h000;
rom[814] = 12'h000;
rom[815] = 12'h000;
rom[816] = 12'h000;
rom[817] = 12'h000;
rom[818] = 12'h000;
rom[819] = 12'h000;
rom[820] = 12'h000;
rom[821] = 12'h000;
rom[822] = 12'h000;
rom[823] = 12'h000;
rom[824] = 12'h00f;
rom[825] = 12'h00f;
rom[826] = 12'h00f;
rom[827] = 12'h00f;
rom[828] = 12'h00f;
rom[829] = 12'h00f;
rom[830] = 12'h000;
rom[831] = 12'h000;
rom[832] = 12'h000;
rom[833] = 12'h000;
rom[834] = 12'h007;
rom[835] = 12'h007;
rom[836] = 12'h000;
rom[837] = 12'h000;
rom[838] = 12'h007;
rom[839] = 12'h007;
rom[840] = 12'h000;
rom[841] = 12'h000;
rom[842] = 12'h000;
rom[843] = 12'h000;
rom[844] = 12'h000;
rom[845] = 12'h000;
rom[846] = 12'h000;
rom[847] = 12'h000;
rom[848] = 12'h000;
rom[849] = 12'h000;
rom[850] = 12'h00f;
rom[851] = 12'h00f;
rom[852] = 12'h00f;
rom[853] = 12'h00f;
rom[854] = 12'h00f;
rom[855] = 12'h00f;
rom[856] = 12'h000;
rom[857] = 12'h000;
rom[858] = 12'h000;
rom[859] = 12'h000;
rom[860] = 12'h007;
rom[861] = 12'h007;
rom[862] = 12'h000;
rom[863] = 12'h000;
rom[864] = 12'h007;
rom[865] = 12'h007;
rom[866] = 12'h000;
rom[867] = 12'h000;
rom[868] = 12'h000;
rom[869] = 12'h000;
rom[870] = 12'h000;
rom[871] = 12'h000;
rom[872] = 12'h000;
rom[873] = 12'h000;
rom[874] = 12'h000;
rom[875] = 12'h000;
rom[876] = 12'h00f;
rom[877] = 12'h00f;
rom[878] = 12'h00f;
rom[879] = 12'h00f;
rom[880] = 12'h00f;
rom[881] = 12'h00f;
rom[882] = 12'h000;
rom[883] = 12'h000;
rom[884] = 12'h000;
rom[885] = 12'h000;
rom[886] = 12'h000;
rom[887] = 12'h000;
rom[888] = 12'h007;
rom[889] = 12'h007;
rom[890] = 12'h000;
rom[891] = 12'h000;
rom[892] = 12'h000;
rom[893] = 12'h000;
rom[894] = 12'h000;
rom[895] = 12'h000;
rom[896] = 12'h000;
rom[897] = 12'h000;
rom[898] = 12'h000;
rom[899] = 12'h000;
rom[900] = 12'h000;
rom[901] = 12'h000;
rom[902] = 12'h00f;
rom[903] = 12'h00f;
rom[904] = 12'h00f;
rom[905] = 12'h00f;
rom[906] = 12'h00f;
rom[907] = 12'h00f;
rom[908] = 12'h000;
rom[909] = 12'h000;
rom[910] = 12'h000;
rom[911] = 12'h000;
rom[912] = 12'h000;
rom[913] = 12'h000;
rom[914] = 12'h007;
rom[915] = 12'h007;
rom[916] = 12'h000;
rom[917] = 12'h000;
rom[918] = 12'h000;
rom[919] = 12'h000;
rom[920] = 12'h000;
rom[921] = 12'h000;
rom[922] = 12'h000;
rom[923] = 12'h000;
rom[924] = 12'h000;
rom[925] = 12'h000;
rom[926] = 12'h000;
rom[927] = 12'h000;
rom[928] = 12'h00f;
rom[929] = 12'h00f;
rom[930] = 12'h00f;
rom[931] = 12'h00f;
rom[932] = 12'h00f;
rom[933] = 12'h00f;
rom[934] = 12'h000;
rom[935] = 12'h000;
rom[936] = 12'h000;
rom[937] = 12'h000;
rom[938] = 12'h007;
rom[939] = 12'h007;
rom[940] = 12'h000;
rom[941] = 12'h000;
rom[942] = 12'h007;
rom[943] = 12'h007;
rom[944] = 12'h000;
rom[945] = 12'h000;
rom[946] = 12'h000;
rom[947] = 12'h000;
rom[948] = 12'h000;
rom[949] = 12'h000;
rom[950] = 12'h000;
rom[951] = 12'h000;
rom[952] = 12'h000;
rom[953] = 12'h000;
rom[954] = 12'h00f;
rom[955] = 12'h00f;
rom[956] = 12'h00f;
rom[957] = 12'h00f;
rom[958] = 12'h00f;
rom[959] = 12'h00f;
rom[960] = 12'h000;
rom[961] = 12'h000;
rom[962] = 12'h000;
rom[963] = 12'h000;
rom[964] = 12'h007;
rom[965] = 12'h007;
rom[966] = 12'h000;
rom[967] = 12'h000;
rom[968] = 12'h007;
rom[969] = 12'h007;
rom[970] = 12'h000;
rom[971] = 12'h000;
rom[972] = 12'h000;
rom[973] = 12'h000;
rom[974] = 12'h000;
rom[975] = 12'h000;
rom[976] = 12'h000;
rom[977] = 12'h000;
rom[978] = 12'h000;
rom[979] = 12'h000;
rom[980] = 12'h00f;
rom[981] = 12'h00f;
rom[982] = 12'h00f;
rom[983] = 12'h00f;
rom[984] = 12'h00f;
rom[985] = 12'h00f;
rom[986] = 12'h000;
rom[987] = 12'h000;
rom[988] = 12'h000;
rom[989] = 12'h000;
rom[990] = 12'h000;
rom[991] = 12'h000;
rom[992] = 12'h007;
rom[993] = 12'h007;
rom[994] = 12'h000;
rom[995] = 12'h000;
rom[996] = 12'h00f;
rom[997] = 12'h00f;
rom[998] = 12'h00f;
rom[999] = 12'h00f;
rom[1000] = 12'h00f;
rom[1001] = 12'h00f;
rom[1002] = 12'h00f;
rom[1003] = 12'h00f;
rom[1004] = 12'h00f;
rom[1005] = 12'h00f;
rom[1006] = 12'h000;
rom[1007] = 12'h000;
rom[1008] = 12'h00f;
rom[1009] = 12'h00f;
rom[1010] = 12'h00f;
rom[1011] = 12'h00f;
rom[1012] = 12'h000;
rom[1013] = 12'h000;
rom[1014] = 12'h000;
rom[1015] = 12'h000;
rom[1016] = 12'h000;
rom[1017] = 12'h000;
rom[1018] = 12'h007;
rom[1019] = 12'h007;
rom[1020] = 12'h000;
rom[1021] = 12'h000;
rom[1022] = 12'h00f;
rom[1023] = 12'h00f;
rom[1024] = 12'h00f;
rom[1025] = 12'h00f;
rom[1026] = 12'h00f;
rom[1027] = 12'h00f;
rom[1028] = 12'h00f;
rom[1029] = 12'h00f;
rom[1030] = 12'h00f;
rom[1031] = 12'h00f;
rom[1032] = 12'h000;
rom[1033] = 12'h000;
rom[1034] = 12'h00f;
rom[1035] = 12'h00f;
rom[1036] = 12'h00f;
rom[1037] = 12'h00f;
rom[1038] = 12'h000;
rom[1039] = 12'h000;
rom[1040] = 12'h000;
rom[1041] = 12'h000;
rom[1042] = 12'h007;
rom[1043] = 12'h007;
rom[1044] = 12'h000;
rom[1045] = 12'h000;
rom[1046] = 12'h00f;
rom[1047] = 12'h00f;
rom[1048] = 12'h00f;
rom[1049] = 12'h00f;
rom[1050] = 12'h00f;
rom[1051] = 12'h00f;
rom[1052] = 12'h00f;
rom[1053] = 12'h00f;
rom[1054] = 12'h00f;
rom[1055] = 12'h00f;
rom[1056] = 12'h00f;
rom[1057] = 12'h00f;
rom[1058] = 12'h00f;
rom[1059] = 12'h00f;
rom[1060] = 12'h000;
rom[1061] = 12'h000;
rom[1062] = 12'h00f;
rom[1063] = 12'h00f;
rom[1064] = 12'h000;
rom[1065] = 12'h000;
rom[1066] = 12'h000;
rom[1067] = 12'h000;
rom[1068] = 12'h007;
rom[1069] = 12'h007;
rom[1070] = 12'h000;
rom[1071] = 12'h000;
rom[1072] = 12'h00f;
rom[1073] = 12'h00f;
rom[1074] = 12'h00f;
rom[1075] = 12'h00f;
rom[1076] = 12'h00f;
rom[1077] = 12'h00f;
rom[1078] = 12'h00f;
rom[1079] = 12'h00f;
rom[1080] = 12'h00f;
rom[1081] = 12'h00f;
rom[1082] = 12'h00f;
rom[1083] = 12'h00f;
rom[1084] = 12'h00f;
rom[1085] = 12'h00f;
rom[1086] = 12'h000;
rom[1087] = 12'h000;
rom[1088] = 12'h00f;
rom[1089] = 12'h00f;
rom[1090] = 12'h000;
rom[1091] = 12'h000;
rom[1092] = 12'h000;
rom[1093] = 12'h000;
rom[1094] = 12'h000;
rom[1095] = 12'h000;
rom[1096] = 12'h00f;
rom[1097] = 12'h00f;
rom[1098] = 12'h00f;
rom[1099] = 12'h00f;
rom[1100] = 12'h00f;
rom[1101] = 12'h00f;
rom[1102] = 12'h00f;
rom[1103] = 12'h00f;
rom[1104] = 12'h00f;
rom[1105] = 12'h00f;
rom[1106] = 12'h00f;
rom[1107] = 12'h00f;
rom[1108] = 12'h00f;
rom[1109] = 12'h00f;
rom[1110] = 12'h00f;
rom[1111] = 12'h00f;
rom[1112] = 12'h00f;
rom[1113] = 12'h00f;
rom[1114] = 12'h000;
rom[1115] = 12'h000;
rom[1116] = 12'h000;
rom[1117] = 12'h000;
rom[1118] = 12'h000;
rom[1119] = 12'h000;
rom[1120] = 12'h000;
rom[1121] = 12'h000;
rom[1122] = 12'h00f;
rom[1123] = 12'h00f;
rom[1124] = 12'h00f;
rom[1125] = 12'h00f;
rom[1126] = 12'h00f;
rom[1127] = 12'h00f;
rom[1128] = 12'h00f;
rom[1129] = 12'h00f;
rom[1130] = 12'h00f;
rom[1131] = 12'h00f;
rom[1132] = 12'h00f;
rom[1133] = 12'h00f;
rom[1134] = 12'h00f;
rom[1135] = 12'h00f;
rom[1136] = 12'h00f;
rom[1137] = 12'h00f;
rom[1138] = 12'h00f;
rom[1139] = 12'h00f;
rom[1140] = 12'h000;
rom[1141] = 12'h000;
rom[1142] = 12'h000;
rom[1143] = 12'h000;
rom[1144] = 12'h000;
rom[1145] = 12'h000;
rom[1146] = 12'h000;
rom[1147] = 12'h000;
rom[1148] = 12'h000;
rom[1149] = 12'h000;
rom[1150] = 12'h000;
rom[1151] = 12'h000;
rom[1152] = 12'h000;
rom[1153] = 12'h000;
rom[1154] = 12'h000;
rom[1155] = 12'h000;
rom[1156] = 12'h000;
rom[1157] = 12'h000;
rom[1158] = 12'h000;
rom[1159] = 12'h000;
rom[1160] = 12'h000;
rom[1161] = 12'h000;
rom[1162] = 12'h000;
rom[1163] = 12'h000;
rom[1164] = 12'h000;
rom[1165] = 12'h000;
rom[1166] = 12'h000;
rom[1167] = 12'h000;
rom[1168] = 12'h000;
rom[1169] = 12'h000;
rom[1170] = 12'h000;
rom[1171] = 12'h000;
rom[1172] = 12'h000;
rom[1173] = 12'h000;
rom[1174] = 12'h000;
rom[1175] = 12'h000;
rom[1176] = 12'h000;
rom[1177] = 12'h000;
rom[1178] = 12'h000;
rom[1179] = 12'h000;
rom[1180] = 12'h000;
rom[1181] = 12'h000;
rom[1182] = 12'h000;
rom[1183] = 12'h000;
rom[1184] = 12'h000;
rom[1185] = 12'h000;
rom[1186] = 12'h000;
rom[1187] = 12'h000;
rom[1188] = 12'h000;
rom[1189] = 12'h000;
rom[1190] = 12'h000;
rom[1191] = 12'h000;
rom[1192] = 12'h000;
rom[1193] = 12'h000;
rom[1194] = 12'h000;
rom[1195] = 12'h000;

  end
  endmodule