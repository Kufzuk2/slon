module tile_mine_exp_rom (                       //невскрытая клетка
  input  wire    [10:0]     addr,
  output wire    [11:0]     word
);

  logic [11:0] rom [(1025)];

  assign word = rom[addr];

  initial begin
rom[0] = 12'h777;
rom[1] = 12'h777;
rom[2] = 12'h777;
rom[3] = 12'h777;
rom[4] = 12'h777;
rom[5] = 12'h777;
rom[6] = 12'h777;
rom[7] = 12'h777;
rom[8] = 12'h777;
rom[9] = 12'h777;
rom[10] = 12'h777;
rom[11] = 12'h777;
rom[12] = 12'h777;
rom[13] = 12'h777;
rom[14] = 12'h777;
rom[15] = 12'h777;
rom[16] = 12'h777;
rom[17] = 12'h777;
rom[18] = 12'h777;
rom[19] = 12'h777;
rom[20] = 12'h777;
rom[21] = 12'h777;
rom[22] = 12'h777;
rom[23] = 12'h777;
rom[24] = 12'h777;
rom[25] = 12'h777;
rom[26] = 12'h777;
rom[27] = 12'h777;
rom[28] = 12'h777;
rom[29] = 12'h777;
rom[30] = 12'h777;
rom[31] = 12'h777;
rom[32] = 12'h777;
rom[33] = 12'h00f;
rom[34] = 12'h00f;
rom[35] = 12'h00f;
rom[36] = 12'h00f;
rom[37] = 12'h00f;
rom[38] = 12'h00f;
rom[39] = 12'h00f;
rom[40] = 12'h00f;
rom[41] = 12'h00f;
rom[42] = 12'h00f;
rom[43] = 12'h00f;
rom[44] = 12'h00f;
rom[45] = 12'h00f;
rom[46] = 12'h00f;
rom[47] = 12'h00f;
rom[48] = 12'h00f;
rom[49] = 12'h00f;
rom[50] = 12'h00f;
rom[51] = 12'h00f;
rom[52] = 12'h00f;
rom[53] = 12'h00f;
rom[54] = 12'h00f;
rom[55] = 12'h00f;
rom[56] = 12'h00f;
rom[57] = 12'h00f;
rom[58] = 12'h00f;
rom[59] = 12'h00f;
rom[60] = 12'h00f;
rom[61] = 12'h00f;
rom[62] = 12'h00f;
rom[63] = 12'h777;
rom[64] = 12'h777;
rom[65] = 12'h00f;
rom[66] = 12'h00f;
rom[67] = 12'h00f;
rom[68] = 12'h00f;
rom[69] = 12'h00f;
rom[70] = 12'h00f;
rom[71] = 12'h00f;
rom[72] = 12'h00f;
rom[73] = 12'h00f;
rom[74] = 12'h00f;
rom[75] = 12'h00f;
rom[76] = 12'h00f;
rom[77] = 12'h00f;
rom[78] = 12'h00f;
rom[79] = 12'h00f;
rom[80] = 12'h00f;
rom[81] = 12'h00f;
rom[82] = 12'h00f;
rom[83] = 12'h00f;
rom[84] = 12'h00f;
rom[85] = 12'h00f;
rom[86] = 12'h00f;
rom[87] = 12'h00f;
rom[88] = 12'h00f;
rom[89] = 12'h00f;
rom[90] = 12'h00f;
rom[91] = 12'h00f;
rom[92] = 12'h00f;
rom[93] = 12'h00f;
rom[94] = 12'h00f;
rom[95] = 12'h777;
rom[96] = 12'h777;
rom[97] = 12'h00f;
rom[98] = 12'h00f;
rom[99] = 12'h00f;
rom[100] = 12'h00f;
rom[101] = 12'h00f;
rom[102] = 12'h00f;
rom[103] = 12'h00f;
rom[104] = 12'h00f;
rom[105] = 12'h00f;
rom[106] = 12'h00f;
rom[107] = 12'h00f;
rom[108] = 12'h00f;
rom[109] = 12'h00f;
rom[110] = 12'h00f;
rom[111] = 12'h00f;
rom[112] = 12'h00f;
rom[113] = 12'h00f;
rom[114] = 12'h00f;
rom[115] = 12'h00f;
rom[116] = 12'h00f;
rom[117] = 12'h00f;
rom[118] = 12'h00f;
rom[119] = 12'h00f;
rom[120] = 12'h00f;
rom[121] = 12'h00f;
rom[122] = 12'h00f;
rom[123] = 12'h00f;
rom[124] = 12'h00f;
rom[125] = 12'h00f;
rom[126] = 12'h00f;
rom[127] = 12'h777;
rom[128] = 12'h777;
rom[129] = 12'h00f;
rom[130] = 12'h00f;
rom[131] = 12'h00f;
rom[132] = 12'h00f;
rom[133] = 12'h00f;
rom[134] = 12'h00f;
rom[135] = 12'h00f;
rom[136] = 12'h00f;
rom[137] = 12'h00f;
rom[138] = 12'h00f;
rom[139] = 12'h00f;
rom[140] = 12'h00f;
rom[141] = 12'h00f;
rom[142] = 12'h00f;
rom[143] = 12'h00f;
rom[144] = 12'h00f;
rom[145] = 12'h00f;
rom[146] = 12'h00f;
rom[147] = 12'h00f;
rom[148] = 12'h00f;
rom[149] = 12'h00f;
rom[150] = 12'h00f;
rom[151] = 12'h00f;
rom[152] = 12'h00f;
rom[153] = 12'h00f;
rom[154] = 12'h00f;
rom[155] = 12'h00f;
rom[156] = 12'h00f;
rom[157] = 12'h00f;
rom[158] = 12'h00f;
rom[159] = 12'h777;
rom[160] = 12'h777;
rom[161] = 12'h00f;
rom[162] = 12'h00f;
rom[163] = 12'h00f;
rom[164] = 12'h00f;
rom[165] = 12'h00f;
rom[166] = 12'h00f;
rom[167] = 12'h00f;
rom[168] = 12'h00f;
rom[169] = 12'h00f;
rom[170] = 12'h00f;
rom[171] = 12'h00f;
rom[172] = 12'h00f;
rom[173] = 12'h00f;
rom[174] = 12'h00f;
rom[175] = 12'h00f;
rom[176] = 12'h00f;
rom[177] = 12'h00f;
rom[178] = 12'h00f;
rom[179] = 12'h00f;
rom[180] = 12'h00f;
rom[181] = 12'h00f;
rom[182] = 12'h00f;
rom[183] = 12'h00f;
rom[184] = 12'h00f;
rom[185] = 12'h00f;
rom[186] = 12'h00f;
rom[187] = 12'h00f;
rom[188] = 12'h00f;
rom[189] = 12'h00f;
rom[190] = 12'h00f;
rom[191] = 12'h777;
rom[192] = 12'h777;
rom[193] = 12'h00f;
rom[194] = 12'h00f;
rom[195] = 12'h00f;
rom[196] = 12'h00f;
rom[197] = 12'h00f;
rom[198] = 12'h00f;
rom[199] = 12'h00f;
rom[200] = 12'h00f;
rom[201] = 12'h00f;
rom[202] = 12'h00f;
rom[203] = 12'h00f;
rom[204] = 12'h00f;
rom[205] = 12'h00f;
rom[206] = 12'h00f;
rom[207] = 12'h00f;
rom[208] = 12'h00f;
rom[209] = 12'h00f;
rom[210] = 12'h00f;
rom[211] = 12'h00f;
rom[212] = 12'h00f;
rom[213] = 12'h00f;
rom[214] = 12'h00f;
rom[215] = 12'h00f;
rom[216] = 12'h00f;
rom[217] = 12'h00f;
rom[218] = 12'h00f;
rom[219] = 12'h00f;
rom[220] = 12'h00f;
rom[221] = 12'h00f;
rom[222] = 12'h00f;
rom[223] = 12'h777;
rom[224] = 12'h777;
rom[225] = 12'h00f;
rom[226] = 12'h00f;
rom[227] = 12'h00f;
rom[228] = 12'h00f;
rom[229] = 12'h00f;
rom[230] = 12'h00f;
rom[231] = 12'h00f;
rom[232] = 12'h00f;
rom[233] = 12'h00f;
rom[234] = 12'h00f;
rom[235] = 12'h00f;
rom[236] = 12'h00f;
rom[237] = 12'h00f;
rom[238] = 12'h00f;
rom[239] = 12'h00f;
rom[240] = 12'h00f;
rom[241] = 12'h00f;
rom[242] = 12'h00f;
rom[243] = 12'h00f;
rom[244] = 12'h00f;
rom[245] = 12'h00f;
rom[246] = 12'h00f;
rom[247] = 12'h00f;
rom[248] = 12'h00f;
rom[249] = 12'h00f;
rom[250] = 12'h00f;
rom[251] = 12'h00f;
rom[252] = 12'h00f;
rom[253] = 12'h00f;
rom[254] = 12'h00f;
rom[255] = 12'h777;
rom[256] = 12'h777;
rom[257] = 12'h00f;
rom[258] = 12'h00f;
rom[259] = 12'h00f;
rom[260] = 12'h00f;
rom[261] = 12'h00f;
rom[262] = 12'h00f;
rom[263] = 12'h00f;
rom[264] = 12'h00f;
rom[265] = 12'h00f;
rom[266] = 12'h00f;
rom[267] = 12'h00f;
rom[268] = 12'h00f;
rom[269] = 12'h00f;
rom[270] = 12'h00f;
rom[271] = 12'h000;
rom[272] = 12'h000;
rom[273] = 12'h00f;
rom[274] = 12'h00f;
rom[275] = 12'h00f;
rom[276] = 12'h00f;
rom[277] = 12'h00f;
rom[278] = 12'h00f;
rom[279] = 12'h00f;
rom[280] = 12'h00f;
rom[281] = 12'h00f;
rom[282] = 12'h00f;
rom[283] = 12'h00f;
rom[284] = 12'h00f;
rom[285] = 12'h00f;
rom[286] = 12'h00f;
rom[287] = 12'h777;
rom[288] = 12'h777;
rom[289] = 12'h00f;
rom[290] = 12'h00f;
rom[291] = 12'h00f;
rom[292] = 12'h00f;
rom[293] = 12'h00f;
rom[294] = 12'h00f;
rom[295] = 12'h00f;
rom[296] = 12'h00f;
rom[297] = 12'h00f;
rom[298] = 12'h00f;
rom[299] = 12'h00f;
rom[300] = 12'h00f;
rom[301] = 12'h00f;
rom[302] = 12'h00f;
rom[303] = 12'h000;
rom[304] = 12'h000;
rom[305] = 12'h00f;
rom[306] = 12'h00f;
rom[307] = 12'h00f;
rom[308] = 12'h00f;
rom[309] = 12'h00f;
rom[310] = 12'h00f;
rom[311] = 12'h00f;
rom[312] = 12'h00f;
rom[313] = 12'h00f;
rom[314] = 12'h00f;
rom[315] = 12'h00f;
rom[316] = 12'h00f;
rom[317] = 12'h00f;
rom[318] = 12'h00f;
rom[319] = 12'h777;
rom[320] = 12'h777;
rom[321] = 12'h00f;
rom[322] = 12'h00f;
rom[323] = 12'h00f;
rom[324] = 12'h00f;
rom[325] = 12'h00f;
rom[326] = 12'h00f;
rom[327] = 12'h00f;
rom[328] = 12'h00f;
rom[329] = 12'h00f;
rom[330] = 12'h000;
rom[331] = 12'h000;
rom[332] = 12'h00f;
rom[333] = 12'h000;
rom[334] = 12'h000;
rom[335] = 12'h000;
rom[336] = 12'h000;
rom[337] = 12'h000;
rom[338] = 12'h000;
rom[339] = 12'h00f;
rom[340] = 12'h000;
rom[341] = 12'h000;
rom[342] = 12'h00f;
rom[343] = 12'h00f;
rom[344] = 12'h00f;
rom[345] = 12'h00f;
rom[346] = 12'h00f;
rom[347] = 12'h00f;
rom[348] = 12'h00f;
rom[349] = 12'h00f;
rom[350] = 12'h00f;
rom[351] = 12'h777;
rom[352] = 12'h777;
rom[353] = 12'h00f;
rom[354] = 12'h00f;
rom[355] = 12'h00f;
rom[356] = 12'h00f;
rom[357] = 12'h00f;
rom[358] = 12'h00f;
rom[359] = 12'h00f;
rom[360] = 12'h00f;
rom[361] = 12'h00f;
rom[362] = 12'h000;
rom[363] = 12'h000;
rom[364] = 12'h00f;
rom[365] = 12'h000;
rom[366] = 12'h000;
rom[367] = 12'h000;
rom[368] = 12'h000;
rom[369] = 12'h000;
rom[370] = 12'h000;
rom[371] = 12'h00f;
rom[372] = 12'h000;
rom[373] = 12'h000;
rom[374] = 12'h00f;
rom[375] = 12'h00f;
rom[376] = 12'h00f;
rom[377] = 12'h00f;
rom[378] = 12'h00f;
rom[379] = 12'h00f;
rom[380] = 12'h00f;
rom[381] = 12'h00f;
rom[382] = 12'h00f;
rom[383] = 12'h777;
rom[384] = 12'h777;
rom[385] = 12'h00f;
rom[386] = 12'h00f;
rom[387] = 12'h00f;
rom[388] = 12'h00f;
rom[389] = 12'h00f;
rom[390] = 12'h00f;
rom[391] = 12'h00f;
rom[392] = 12'h00f;
rom[393] = 12'h00f;
rom[394] = 12'h00f;
rom[395] = 12'h00f;
rom[396] = 12'h000;
rom[397] = 12'h000;
rom[398] = 12'h000;
rom[399] = 12'h000;
rom[400] = 12'h000;
rom[401] = 12'h000;
rom[402] = 12'h000;
rom[403] = 12'h000;
rom[404] = 12'h00f;
rom[405] = 12'h00f;
rom[406] = 12'h00f;
rom[407] = 12'h00f;
rom[408] = 12'h00f;
rom[409] = 12'h00f;
rom[410] = 12'h00f;
rom[411] = 12'h00f;
rom[412] = 12'h00f;
rom[413] = 12'h00f;
rom[414] = 12'h00f;
rom[415] = 12'h777;
rom[416] = 12'h777;
rom[417] = 12'h00f;
rom[418] = 12'h00f;
rom[419] = 12'h00f;
rom[420] = 12'h00f;
rom[421] = 12'h00f;
rom[422] = 12'h00f;
rom[423] = 12'h00f;
rom[424] = 12'h00f;
rom[425] = 12'h00f;
rom[426] = 12'h000;
rom[427] = 12'h000;
rom[428] = 12'h000;
rom[429] = 12'hfff;
rom[430] = 12'hfff;
rom[431] = 12'h000;
rom[432] = 12'h000;
rom[433] = 12'h000;
rom[434] = 12'h000;
rom[435] = 12'h000;
rom[436] = 12'h000;
rom[437] = 12'h000;
rom[438] = 12'h00f;
rom[439] = 12'h00f;
rom[440] = 12'h00f;
rom[441] = 12'h00f;
rom[442] = 12'h00f;
rom[443] = 12'h00f;
rom[444] = 12'h00f;
rom[445] = 12'h00f;
rom[446] = 12'h00f;
rom[447] = 12'h777;
rom[448] = 12'h777;
rom[449] = 12'h00f;
rom[450] = 12'h00f;
rom[451] = 12'h00f;
rom[452] = 12'h00f;
rom[453] = 12'h00f;
rom[454] = 12'h00f;
rom[455] = 12'h00f;
rom[456] = 12'h00f;
rom[457] = 12'h00f;
rom[458] = 12'h000;
rom[459] = 12'h000;
rom[460] = 12'h000;
rom[461] = 12'hfff;
rom[462] = 12'hfff;
rom[463] = 12'h000;
rom[464] = 12'h000;
rom[465] = 12'h000;
rom[466] = 12'h000;
rom[467] = 12'h000;
rom[468] = 12'h000;
rom[469] = 12'h000;
rom[470] = 12'h00f;
rom[471] = 12'h00f;
rom[472] = 12'h00f;
rom[473] = 12'h00f;
rom[474] = 12'h00f;
rom[475] = 12'h00f;
rom[476] = 12'h00f;
rom[477] = 12'h00f;
rom[478] = 12'h00f;
rom[479] = 12'h777;
rom[480] = 12'h777;
rom[481] = 12'h00f;
rom[482] = 12'h00f;
rom[483] = 12'h00f;
rom[484] = 12'h00f;
rom[485] = 12'h00f;
rom[486] = 12'h00f;
rom[487] = 12'h00f;
rom[488] = 12'h000;
rom[489] = 12'h000;
rom[490] = 12'h000;
rom[491] = 12'h000;
rom[492] = 12'h000;
rom[493] = 12'h000;
rom[494] = 12'h000;
rom[495] = 12'h000;
rom[496] = 12'h000;
rom[497] = 12'h000;
rom[498] = 12'h000;
rom[499] = 12'h000;
rom[500] = 12'h000;
rom[501] = 12'h000;
rom[502] = 12'h000;
rom[503] = 12'h000;
rom[504] = 12'h00f;
rom[505] = 12'h00f;
rom[506] = 12'h00f;
rom[507] = 12'h00f;
rom[508] = 12'h00f;
rom[509] = 12'h00f;
rom[510] = 12'h00f;
rom[511] = 12'h777;
rom[512] = 12'h777;
rom[513] = 12'h00f;
rom[514] = 12'h00f;
rom[515] = 12'h00f;
rom[516] = 12'h00f;
rom[517] = 12'h00f;
rom[518] = 12'h00f;
rom[519] = 12'h00f;
rom[520] = 12'h000;
rom[521] = 12'h000;
rom[522] = 12'h000;
rom[523] = 12'h000;
rom[524] = 12'h000;
rom[525] = 12'h000;
rom[526] = 12'h000;
rom[527] = 12'h000;
rom[528] = 12'h000;
rom[529] = 12'h000;
rom[530] = 12'h000;
rom[531] = 12'h000;
rom[532] = 12'h000;
rom[533] = 12'h000;
rom[534] = 12'h000;
rom[535] = 12'h000;
rom[536] = 12'h00f;
rom[537] = 12'h00f;
rom[538] = 12'h00f;
rom[539] = 12'h00f;
rom[540] = 12'h00f;
rom[541] = 12'h00f;
rom[542] = 12'h00f;
rom[543] = 12'h777;
rom[544] = 12'h777;
rom[545] = 12'h00f;
rom[546] = 12'h00f;
rom[547] = 12'h00f;
rom[548] = 12'h00f;
rom[549] = 12'h00f;
rom[550] = 12'h00f;
rom[551] = 12'h00f;
rom[552] = 12'h00f;
rom[553] = 12'h00f;
rom[554] = 12'h000;
rom[555] = 12'h000;
rom[556] = 12'h000;
rom[557] = 12'h000;
rom[558] = 12'h000;
rom[559] = 12'h000;
rom[560] = 12'h000;
rom[561] = 12'h000;
rom[562] = 12'h000;
rom[563] = 12'h000;
rom[564] = 12'h000;
rom[565] = 12'h000;
rom[566] = 12'h00f;
rom[567] = 12'h00f;
rom[568] = 12'h00f;
rom[569] = 12'h00f;
rom[570] = 12'h00f;
rom[571] = 12'h00f;
rom[572] = 12'h00f;
rom[573] = 12'h00f;
rom[574] = 12'h00f;
rom[575] = 12'h777;
rom[576] = 12'h777;
rom[577] = 12'h00f;
rom[578] = 12'h00f;
rom[579] = 12'h00f;
rom[580] = 12'h00f;
rom[581] = 12'h00f;
rom[582] = 12'h00f;
rom[583] = 12'h00f;
rom[584] = 12'h00f;
rom[585] = 12'h00f;
rom[586] = 12'h000;
rom[587] = 12'h000;
rom[588] = 12'h000;
rom[589] = 12'h000;
rom[590] = 12'h000;
rom[591] = 12'h000;
rom[592] = 12'h000;
rom[593] = 12'h000;
rom[594] = 12'h000;
rom[595] = 12'h000;
rom[596] = 12'h000;
rom[597] = 12'h000;
rom[598] = 12'h00f;
rom[599] = 12'h00f;
rom[600] = 12'h00f;
rom[601] = 12'h00f;
rom[602] = 12'h00f;
rom[603] = 12'h00f;
rom[604] = 12'h00f;
rom[605] = 12'h00f;
rom[606] = 12'h00f;
rom[607] = 12'h777;
rom[608] = 12'h777;
rom[609] = 12'h00f;
rom[610] = 12'h00f;
rom[611] = 12'h00f;
rom[612] = 12'h00f;
rom[613] = 12'h00f;
rom[614] = 12'h00f;
rom[615] = 12'h00f;
rom[616] = 12'h00f;
rom[617] = 12'h00f;
rom[618] = 12'h00f;
rom[619] = 12'h00f;
rom[620] = 12'h000;
rom[621] = 12'h000;
rom[622] = 12'h000;
rom[623] = 12'h000;
rom[624] = 12'h000;
rom[625] = 12'h000;
rom[626] = 12'h000;
rom[627] = 12'h000;
rom[628] = 12'h00f;
rom[629] = 12'h00f;
rom[630] = 12'h00f;
rom[631] = 12'h00f;
rom[632] = 12'h00f;
rom[633] = 12'h00f;
rom[634] = 12'h00f;
rom[635] = 12'h00f;
rom[636] = 12'h00f;
rom[637] = 12'h00f;
rom[638] = 12'h00f;
rom[639] = 12'h777;
rom[640] = 12'h777;
rom[641] = 12'h00f;
rom[642] = 12'h00f;
rom[643] = 12'h00f;
rom[644] = 12'h00f;
rom[645] = 12'h00f;
rom[646] = 12'h00f;
rom[647] = 12'h00f;
rom[648] = 12'h00f;
rom[649] = 12'h00f;
rom[650] = 12'h000;
rom[651] = 12'h000;
rom[652] = 12'h00f;
rom[653] = 12'h000;
rom[654] = 12'h000;
rom[655] = 12'h000;
rom[656] = 12'h000;
rom[657] = 12'h000;
rom[658] = 12'h000;
rom[659] = 12'h00f;
rom[660] = 12'h000;
rom[661] = 12'h000;
rom[662] = 12'h00f;
rom[663] = 12'h00f;
rom[664] = 12'h00f;
rom[665] = 12'h00f;
rom[666] = 12'h00f;
rom[667] = 12'h00f;
rom[668] = 12'h00f;
rom[669] = 12'h00f;
rom[670] = 12'h00f;
rom[671] = 12'h777;
rom[672] = 12'h777;
rom[673] = 12'h00f;
rom[674] = 12'h00f;
rom[675] = 12'h00f;
rom[676] = 12'h00f;
rom[677] = 12'h00f;
rom[678] = 12'h00f;
rom[679] = 12'h00f;
rom[680] = 12'h00f;
rom[681] = 12'h00f;
rom[682] = 12'h000;
rom[683] = 12'h000;
rom[684] = 12'h00f;
rom[685] = 12'h000;
rom[686] = 12'h000;
rom[687] = 12'h000;
rom[688] = 12'h000;
rom[689] = 12'h000;
rom[690] = 12'h000;
rom[691] = 12'h00f;
rom[692] = 12'h000;
rom[693] = 12'h000;
rom[694] = 12'h00f;
rom[695] = 12'h00f;
rom[696] = 12'h00f;
rom[697] = 12'h00f;
rom[698] = 12'h00f;
rom[699] = 12'h00f;
rom[700] = 12'h00f;
rom[701] = 12'h00f;
rom[702] = 12'h00f;
rom[703] = 12'h777;
rom[704] = 12'h777;
rom[705] = 12'h00f;
rom[706] = 12'h00f;
rom[707] = 12'h00f;
rom[708] = 12'h00f;
rom[709] = 12'h00f;
rom[710] = 12'h00f;
rom[711] = 12'h00f;
rom[712] = 12'h00f;
rom[713] = 12'h00f;
rom[714] = 12'h00f;
rom[715] = 12'h00f;
rom[716] = 12'h00f;
rom[717] = 12'h00f;
rom[718] = 12'h00f;
rom[719] = 12'h000;
rom[720] = 12'h000;
rom[721] = 12'h00f;
rom[722] = 12'h00f;
rom[723] = 12'h00f;
rom[724] = 12'h00f;
rom[725] = 12'h00f;
rom[726] = 12'h00f;
rom[727] = 12'h00f;
rom[728] = 12'h00f;
rom[729] = 12'h00f;
rom[730] = 12'h00f;
rom[731] = 12'h00f;
rom[732] = 12'h00f;
rom[733] = 12'h00f;
rom[734] = 12'h00f;
rom[735] = 12'h777;
rom[736] = 12'h777;
rom[737] = 12'h00f;
rom[738] = 12'h00f;
rom[739] = 12'h00f;
rom[740] = 12'h00f;
rom[741] = 12'h00f;
rom[742] = 12'h00f;
rom[743] = 12'h00f;
rom[744] = 12'h00f;
rom[745] = 12'h00f;
rom[746] = 12'h00f;
rom[747] = 12'h00f;
rom[748] = 12'h00f;
rom[749] = 12'h00f;
rom[750] = 12'h00f;
rom[751] = 12'h000;
rom[752] = 12'h000;
rom[753] = 12'h00f;
rom[754] = 12'h00f;
rom[755] = 12'h00f;
rom[756] = 12'h00f;
rom[757] = 12'h00f;
rom[758] = 12'h00f;
rom[759] = 12'h00f;
rom[760] = 12'h00f;
rom[761] = 12'h00f;
rom[762] = 12'h00f;
rom[763] = 12'h00f;
rom[764] = 12'h00f;
rom[765] = 12'h00f;
rom[766] = 12'h00f;
rom[767] = 12'h777;
rom[768] = 12'h777;
rom[769] = 12'h00f;
rom[770] = 12'h00f;
rom[771] = 12'h00f;
rom[772] = 12'h00f;
rom[773] = 12'h00f;
rom[774] = 12'h00f;
rom[775] = 12'h00f;
rom[776] = 12'h00f;
rom[777] = 12'h00f;
rom[778] = 12'h00f;
rom[779] = 12'h00f;
rom[780] = 12'h00f;
rom[781] = 12'h00f;
rom[782] = 12'h00f;
rom[783] = 12'h00f;
rom[784] = 12'h00f;
rom[785] = 12'h00f;
rom[786] = 12'h00f;
rom[787] = 12'h00f;
rom[788] = 12'h00f;
rom[789] = 12'h00f;
rom[790] = 12'h00f;
rom[791] = 12'h00f;
rom[792] = 12'h00f;
rom[793] = 12'h00f;
rom[794] = 12'h00f;
rom[795] = 12'h00f;
rom[796] = 12'h00f;
rom[797] = 12'h00f;
rom[798] = 12'h00f;
rom[799] = 12'h777;
rom[800] = 12'h777;
rom[801] = 12'h00f;
rom[802] = 12'h00f;
rom[803] = 12'h00f;
rom[804] = 12'h00f;
rom[805] = 12'h00f;
rom[806] = 12'h00f;
rom[807] = 12'h00f;
rom[808] = 12'h00f;
rom[809] = 12'h00f;
rom[810] = 12'h00f;
rom[811] = 12'h00f;
rom[812] = 12'h00f;
rom[813] = 12'h00f;
rom[814] = 12'h00f;
rom[815] = 12'h00f;
rom[816] = 12'h00f;
rom[817] = 12'h00f;
rom[818] = 12'h00f;
rom[819] = 12'h00f;
rom[820] = 12'h00f;
rom[821] = 12'h00f;
rom[822] = 12'h00f;
rom[823] = 12'h00f;
rom[824] = 12'h00f;
rom[825] = 12'h00f;
rom[826] = 12'h00f;
rom[827] = 12'h00f;
rom[828] = 12'h00f;
rom[829] = 12'h00f;
rom[830] = 12'h00f;
rom[831] = 12'h777;
rom[832] = 12'h777;
rom[833] = 12'h00f;
rom[834] = 12'h00f;
rom[835] = 12'h00f;
rom[836] = 12'h00f;
rom[837] = 12'h00f;
rom[838] = 12'h00f;
rom[839] = 12'h00f;
rom[840] = 12'h00f;
rom[841] = 12'h00f;
rom[842] = 12'h00f;
rom[843] = 12'h00f;
rom[844] = 12'h00f;
rom[845] = 12'h00f;
rom[846] = 12'h00f;
rom[847] = 12'h00f;
rom[848] = 12'h00f;
rom[849] = 12'h00f;
rom[850] = 12'h00f;
rom[851] = 12'h00f;
rom[852] = 12'h00f;
rom[853] = 12'h00f;
rom[854] = 12'h00f;
rom[855] = 12'h00f;
rom[856] = 12'h00f;
rom[857] = 12'h00f;
rom[858] = 12'h00f;
rom[859] = 12'h00f;
rom[860] = 12'h00f;
rom[861] = 12'h00f;
rom[862] = 12'h00f;
rom[863] = 12'h777;
rom[864] = 12'h777;
rom[865] = 12'h00f;
rom[866] = 12'h00f;
rom[867] = 12'h00f;
rom[868] = 12'h00f;
rom[869] = 12'h00f;
rom[870] = 12'h00f;
rom[871] = 12'h00f;
rom[872] = 12'h00f;
rom[873] = 12'h00f;
rom[874] = 12'h00f;
rom[875] = 12'h00f;
rom[876] = 12'h00f;
rom[877] = 12'h00f;
rom[878] = 12'h00f;
rom[879] = 12'h00f;
rom[880] = 12'h00f;
rom[881] = 12'h00f;
rom[882] = 12'h00f;
rom[883] = 12'h00f;
rom[884] = 12'h00f;
rom[885] = 12'h00f;
rom[886] = 12'h00f;
rom[887] = 12'h00f;
rom[888] = 12'h00f;
rom[889] = 12'h00f;
rom[890] = 12'h00f;
rom[891] = 12'h00f;
rom[892] = 12'h00f;
rom[893] = 12'h00f;
rom[894] = 12'h00f;
rom[895] = 12'h777;
rom[896] = 12'h777;
rom[897] = 12'h00f;
rom[898] = 12'h00f;
rom[899] = 12'h00f;
rom[900] = 12'h00f;
rom[901] = 12'h00f;
rom[902] = 12'h00f;
rom[903] = 12'h00f;
rom[904] = 12'h00f;
rom[905] = 12'h00f;
rom[906] = 12'h00f;
rom[907] = 12'h00f;
rom[908] = 12'h00f;
rom[909] = 12'h00f;
rom[910] = 12'h00f;
rom[911] = 12'h00f;
rom[912] = 12'h00f;
rom[913] = 12'h00f;
rom[914] = 12'h00f;
rom[915] = 12'h00f;
rom[916] = 12'h00f;
rom[917] = 12'h00f;
rom[918] = 12'h00f;
rom[919] = 12'h00f;
rom[920] = 12'h00f;
rom[921] = 12'h00f;
rom[922] = 12'h00f;
rom[923] = 12'h00f;
rom[924] = 12'h00f;
rom[925] = 12'h00f;
rom[926] = 12'h00f;
rom[927] = 12'h777;
rom[928] = 12'h777;
rom[929] = 12'h00f;
rom[930] = 12'h00f;
rom[931] = 12'h00f;
rom[932] = 12'h00f;
rom[933] = 12'h00f;
rom[934] = 12'h00f;
rom[935] = 12'h00f;
rom[936] = 12'h00f;
rom[937] = 12'h00f;
rom[938] = 12'h00f;
rom[939] = 12'h00f;
rom[940] = 12'h00f;
rom[941] = 12'h00f;
rom[942] = 12'h00f;
rom[943] = 12'h00f;
rom[944] = 12'h00f;
rom[945] = 12'h00f;
rom[946] = 12'h00f;
rom[947] = 12'h00f;
rom[948] = 12'h00f;
rom[949] = 12'h00f;
rom[950] = 12'h00f;
rom[951] = 12'h00f;
rom[952] = 12'h00f;
rom[953] = 12'h00f;
rom[954] = 12'h00f;
rom[955] = 12'h00f;
rom[956] = 12'h00f;
rom[957] = 12'h00f;
rom[958] = 12'h00f;
rom[959] = 12'h777;
rom[960] = 12'h777;
rom[961] = 12'h00f;
rom[962] = 12'h00f;
rom[963] = 12'h00f;
rom[964] = 12'h00f;
rom[965] = 12'h00f;
rom[966] = 12'h00f;
rom[967] = 12'h00f;
rom[968] = 12'h00f;
rom[969] = 12'h00f;
rom[970] = 12'h00f;
rom[971] = 12'h00f;
rom[972] = 12'h00f;
rom[973] = 12'h00f;
rom[974] = 12'h00f;
rom[975] = 12'h00f;
rom[976] = 12'h00f;
rom[977] = 12'h00f;
rom[978] = 12'h00f;
rom[979] = 12'h00f;
rom[980] = 12'h00f;
rom[981] = 12'h00f;
rom[982] = 12'h00f;
rom[983] = 12'h00f;
rom[984] = 12'h00f;
rom[985] = 12'h00f;
rom[986] = 12'h00f;
rom[987] = 12'h00f;
rom[988] = 12'h00f;
rom[989] = 12'h00f;
rom[990] = 12'h00f;
rom[991] = 12'h777;
rom[992] = 12'h777;
rom[993] = 12'h777;
rom[994] = 12'h777;
rom[995] = 12'h777;
rom[996] = 12'h777;
rom[997] = 12'h777;
rom[998] = 12'h777;
rom[999] = 12'h777;
rom[1000] = 12'h777;
rom[1001] = 12'h777;
rom[1002] = 12'h777;
rom[1003] = 12'h777;
rom[1004] = 12'h777;
rom[1005] = 12'h777;
rom[1006] = 12'h777;
rom[1007] = 12'h777;
rom[1008] = 12'h777;
rom[1009] = 12'h777;
rom[1010] = 12'h777;
rom[1011] = 12'h777;
rom[1012] = 12'h777;
rom[1013] = 12'h777;
rom[1014] = 12'h777;
rom[1015] = 12'h777;
rom[1016] = 12'h777;
rom[1017] = 12'h777;
rom[1018] = 12'h777;
rom[1019] = 12'h777;
rom[1020] = 12'h777;
rom[1021] = 12'h777;
rom[1022] = 12'h777;
rom[1023] = 12'h777;
  end

endmodule